** Generated for: hspiceD
** Generated on: Dec  6 20:51:35 2016
** Design library name: Project_416
** Design cell name: CBA_16bit
** Design view name: extracted


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20N.m"
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20P.m"

** Library name: Project_416
** Cell name: CBA_16bit
** View name: extracted
m0 n56 n125 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m1 vdd n57 n56 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m2 n65 n135 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m3 vdd n202 n65 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m4 n79 a8 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m5 vdd b8 n79 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m6 n86 b7 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m7 vdd a7 n86 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m8 n94 a9 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m9 vdd b9 n94 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m10 n101 b6 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m11 vdd a6 n101 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m12 n160 a10 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m13 vdd b10 n160 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m14 n167 b5 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m15 vdd a5 n167 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m16 n175 a11 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m17 vdd b11 n175 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m18 n182 b4 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m19 vdd a4 n182 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m20 n197 n53 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m21 vdd n116 n197 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m22 n206 n198 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m23 vdd n128 n206 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m24 n212 n281 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m25 vdd n213 n212 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m26 n221 n291 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m27 vdd n358 n221 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m28 n235 a12 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m29 vdd b12 n235 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m30 n242 b3 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m31 vdd a3 n242 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m32 n250 a13 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m33 vdd b13 n250 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m34 n257 b2 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m35 vdd a2 n257 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m36 n316 a14 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m37 vdd b14 n316 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m38 n323 b1 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m39 vdd a1 n323 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m40 n331 a15 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m41 vdd b15 n331 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m42 n338 b0 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m43 vdd a0 n338 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m44 n353 n209 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m45 vdd n272 n353 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
m46 n361 n354 vdd vdd tsmc20P L=200e-9 W=900e-9 AD=270e-15 AS=450e-15 PD=600e-9 PS=1.9e-6 M=1
m47 vdd n284 n361 vdd tsmc20P L=200e-9 W=900e-9 AD=450e-15 AS=270e-15 PD=1.9e-6 PS=600e-9 M=1
c48 gnd n361 45.59e-18 M=1
c49 gnd n358 153.26e-18 M=1
c50 gnd n357 95.06e-18 M=1
c51 gnd n356 73.72e-18 M=1
c52 gnd n354 157.14e-18 M=1
c53 gnd n353 45.59e-18 M=1
c54 gnd n350 73.72e-18 M=1
c55 gnd n349 67.9e-18 M=1
c56 gnd n348 73.72e-18 M=1
c57 gnd n346 25.22e-18 M=1
c58 gnd n345 73.72e-18 M=1
c59 gnd n344 73.72e-18 M=1
c60 gnd n343 60.14e-18 M=1
c61 gnd n342 73.72e-18 M=1
c62 gnd n340 73.72e-18 M=1
c63 gnd n338 21.34e-18 M=1
c64 gnd n337 54.32e-18 M=1
c65 gnd n335 54.32e-18 M=1
c66 gnd n333 73.72e-18 M=1
c67 gnd n332 25.22e-18 M=1
c68 gnd n331 21.34e-18 M=1
c69 gnd n330 25.22e-18 M=1
c70 gnd n328 120.28e-18 M=1
c71 gnd n327 60.14e-18 M=1
c72 gnd n324 25.22e-18 M=1
c73 gnd n323 21.34e-18 M=1
c74 gnd n322 25.22e-18 M=1
c75 gnd n321 73.72e-18 M=1
c76 gnd n318 67.9e-18 M=1
c77 gnd n317 67.9e-18 M=1
c78 gnd n316 21.34e-18 M=1
c79 gnd n315 73.72e-18 M=1
c80 gnd n313 73.72e-18 M=1
c81 gnd n312 73.72e-18 M=1
c82 gnd n311 60.14e-18 M=1
c83 gnd n310 120.28e-18 M=1
c84 gnd n307 73.72e-18 M=1
c85 gnd n306 73.72e-18 M=1
c86 gnd n305 73.72e-18 M=1
c87 gnd n304 54.32e-18 M=1
c88 gnd n303 54.32e-18 M=1
c89 gnd n299 73.72e-18 M=1
c90 gnd n298 120.28e-18 M=1
c91 gnd n297 60.14e-18 M=1
c92 gnd n296 73.72e-18 M=1
c93 gnd n291 157.14e-18 M=1
c94 gnd n290 67.9e-18 M=1
c95 gnd n289 73.72e-18 M=1
c96 gnd n286 73.72e-18 M=1
c97 gnd n285 67.9e-18 M=1
c98 gnd n284 153.26e-18 M=1
c99 gnd n281 153.26e-18 M=1
c100 gnd n279 73.72e-18 M=1
c101 gnd n278 60.14e-18 M=1
c102 gnd n277 120.28e-18 M=1
c103 gnd n276 73.72e-18 M=1
c104 gnd n272 157.14e-18 M=1
c105 gnd n270 54.32e-18 M=1
c106 gnd n269 54.32e-18 M=1
c107 gnd n268 73.72e-18 M=1
c108 gnd n267 73.72e-18 M=1
c109 gnd n266 73.72e-18 M=1
c110 gnd n264 120.28e-18 M=1
c111 gnd n263 60.14e-18 M=1
c112 gnd n261 73.72e-18 M=1
c113 gnd n260 73.72e-18 M=1
c114 gnd n258 73.72e-18 M=1
c115 gnd n257 21.34e-18 M=1
c116 gnd n256 67.9e-18 M=1
c117 gnd n255 67.9e-18 M=1
c118 gnd n252 73.72e-18 M=1
c119 gnd n251 25.22e-18 M=1
c120 gnd n250 21.34e-18 M=1
c121 gnd n249 25.22e-18 M=1
c122 gnd n247 60.14e-18 M=1
c123 gnd n246 120.28e-18 M=1
c124 gnd n244 25.22e-18 M=1
c125 gnd n242 21.34e-18 M=1
c126 gnd n241 25.22e-18 M=1
c127 gnd n240 73.72e-18 M=1
c128 gnd n238 54.32e-18 M=1
c129 gnd n236 54.32e-18 M=1
c130 gnd n235 21.34e-18 M=1
c131 gnd n234 73.72e-18 M=1
c132 gnd n232 73.72e-18 M=1
c133 gnd n231 60.14e-18 M=1
c134 gnd n230 73.72e-18 M=1
c135 gnd n229 73.72e-18 M=1
c136 gnd n226 73.72e-18 M=1
c137 gnd n225 67.9e-18 M=1
c138 gnd n224 73.72e-18 M=1
c139 gnd n221 45.59e-18 M=1
c140 gnd n220 25.22e-18 M=1
c141 gnd n218 73.72e-18 M=1
c142 gnd n217 95.06e-18 M=1
c143 gnd n215 194e-18 M=1
c144 gnd n213 157.14e-18 M=1
c145 gnd n212 45.59e-18 M=1
c146 gnd n209 153.26e-18 M=1
c147 gnd n206 45.59e-18 M=1
c148 gnd n204 194e-18 M=1
c149 gnd n202 153.26e-18 M=1
c150 gnd n201 95.06e-18 M=1
c151 gnd n200 73.72e-18 M=1
c152 gnd n198 157.14e-18 M=1
c153 gnd n197 45.59e-18 M=1
c154 gnd n194 73.72e-18 M=1
c155 gnd n193 67.9e-18 M=1
c156 gnd n192 73.72e-18 M=1
c157 gnd n190 25.22e-18 M=1
c158 gnd n189 73.72e-18 M=1
c159 gnd n188 73.72e-18 M=1
c160 gnd n187 60.14e-18 M=1
c161 gnd n186 73.72e-18 M=1
c162 gnd n184 73.72e-18 M=1
c163 gnd n182 21.34e-18 M=1
c164 gnd n181 54.32e-18 M=1
c165 gnd n179 54.32e-18 M=1
c166 gnd n177 73.72e-18 M=1
c167 gnd n176 25.22e-18 M=1
c168 gnd n175 21.34e-18 M=1
c169 gnd n174 25.22e-18 M=1
c170 gnd n172 120.28e-18 M=1
c171 gnd n171 60.14e-18 M=1
c172 gnd n168 25.22e-18 M=1
c173 gnd n167 21.34e-18 M=1
c174 gnd n166 25.22e-18 M=1
c175 gnd n165 73.72e-18 M=1
c176 gnd n162 67.9e-18 M=1
c177 gnd n161 67.9e-18 M=1
c178 gnd n160 21.34e-18 M=1
c179 gnd n159 73.72e-18 M=1
c180 gnd n157 73.72e-18 M=1
c181 gnd n156 73.72e-18 M=1
c182 gnd n155 60.14e-18 M=1
c183 gnd n154 120.28e-18 M=1
c184 gnd n151 73.72e-18 M=1
c185 gnd n150 73.72e-18 M=1
c186 gnd n149 73.72e-18 M=1
c187 gnd n148 54.32e-18 M=1
c188 gnd n147 54.32e-18 M=1
c189 gnd n143 73.72e-18 M=1
c190 gnd n142 120.28e-18 M=1
c191 gnd n141 60.14e-18 M=1
c192 gnd n140 73.72e-18 M=1
c193 gnd n135 157.14e-18 M=1
c194 gnd n134 67.9e-18 M=1
c195 gnd n133 73.72e-18 M=1
c196 gnd n130 73.72e-18 M=1
c197 gnd n129 67.9e-18 M=1
c198 gnd n128 153.26e-18 M=1
c199 gnd n125 153.26e-18 M=1
c200 gnd n123 73.72e-18 M=1
c201 gnd n122 60.14e-18 M=1
c202 gnd n121 120.28e-18 M=1
c203 gnd n120 73.72e-18 M=1
c204 gnd n116 157.14e-18 M=1
c205 gnd n114 54.32e-18 M=1
c206 gnd n113 54.32e-18 M=1
c207 gnd n112 73.72e-18 M=1
c208 gnd n111 73.72e-18 M=1
c209 gnd n110 73.72e-18 M=1
c210 gnd n108 120.28e-18 M=1
c211 gnd n107 60.14e-18 M=1
c212 gnd n105 73.72e-18 M=1
c213 gnd n104 73.72e-18 M=1
c214 gnd n102 73.72e-18 M=1
c215 gnd n101 21.34e-18 M=1
c216 gnd n100 67.9e-18 M=1
c217 gnd n99 67.9e-18 M=1
c218 gnd n96 73.72e-18 M=1
c219 gnd n95 25.22e-18 M=1
c220 gnd n94 21.34e-18 M=1
c221 gnd n93 25.22e-18 M=1
c222 gnd n91 60.14e-18 M=1
c223 gnd n90 120.28e-18 M=1
c224 gnd n88 25.22e-18 M=1
c225 gnd n86 21.34e-18 M=1
c226 gnd n85 25.22e-18 M=1
c227 gnd n84 73.72e-18 M=1
c228 gnd n82 54.32e-18 M=1
c229 gnd n80 54.32e-18 M=1
c230 gnd n79 21.34e-18 M=1
c231 gnd n78 73.72e-18 M=1
c232 gnd n76 73.72e-18 M=1
c233 gnd n75 60.14e-18 M=1
c234 gnd n74 73.72e-18 M=1
c235 gnd n73 73.72e-18 M=1
c236 gnd n70 73.72e-18 M=1
c237 gnd n69 67.9e-18 M=1
c238 gnd n68 73.72e-18 M=1
c239 gnd n65 45.59e-18 M=1
c240 gnd n64 25.22e-18 M=1
c241 gnd n62 73.72e-18 M=1
c242 gnd n61 95.06e-18 M=1
c243 gnd n59 194e-18 M=1
c244 gnd n57 157.14e-18 M=1
c245 gnd n56 45.59e-18 M=1
c246 gnd n53 153.26e-18 M=1
c247 gnd a9 131.92e-18 M=1
c248 gnd a8 124.16e-18 M=1
c249 gnd a7 131.92e-18 M=1
c250 gnd a6 124.16e-18 M=1
c251 gnd a5 131.92e-18 M=1
c252 gnd a4 124.16e-18 M=1
c253 gnd a3 131.92e-18 M=1
c254 gnd a2 124.16e-18 M=1
c255 gnd a1 131.92e-18 M=1
c256 gnd a0 124.16e-18 M=1
c257 gnd b15 124.16e-18 M=1
c258 gnd b14 131.92e-18 M=1
c259 gnd b13 124.16e-18 M=1
c260 gnd b12 131.92e-18 M=1
c261 gnd b11 124.16e-18 M=1
c262 gnd b10 131.92e-18 M=1
c263 a15 gnd 131.92e-18 M=1
c264 a14 gnd 124.16e-18 M=1
c265 a13 gnd 131.92e-18 M=1
c266 a12 gnd 124.16e-18 M=1
c267 a11 gnd 131.92e-18 M=1
c268 a10 gnd 124.16e-18 M=1
c269 cin gnd 194e-18 M=1
c270 b9 gnd 124.16e-18 M=1
c271 b8 gnd 131.92e-18 M=1
c272 b7 gnd 124.16e-18 M=1
c273 b6 gnd 131.92e-18 M=1
c274 b5 gnd 124.16e-18 M=1
c275 b4 gnd 131.92e-18 M=1
c276 b3 gnd 124.16e-18 M=1
c277 b2 gnd 131.92e-18 M=1
c278 b1 gnd 124.16e-18 M=1
c279 b0 gnd 131.92e-18 M=1
c280 vdd n358 89.24e-18 M=1
c281 vdd n357 50.44e-18 M=1
c282 vdd n354 77.6e-18 M=1
c283 vdd n346 23.28e-18 M=1
c284 vdd n338 27.16e-18 M=1
c285 vdd n337 21.34e-18 M=1
c286 vdd n335 21.34e-18 M=1
c287 vdd n332 23.28e-18 M=1
c288 vdd n331 27.16e-18 M=1
c289 vdd n330 23.28e-18 M=1
c290 vdd n328 73.72e-18 M=1
c291 vdd n324 23.28e-18 M=1
c292 vdd n323 27.16e-18 M=1
c293 vdd n322 23.28e-18 M=1
c294 vdd n316 27.16e-18 M=1
c295 vdd n310 73.72e-18 M=1
c296 vdd n304 21.34e-18 M=1
c297 vdd n303 21.34e-18 M=1
c298 vdd n298 73.72e-18 M=1
c299 vdd n291 77.6e-18 M=1
c300 vdd n284 89.24e-18 M=1
c301 vdd n281 89.24e-18 M=1
c302 vdd n277 73.72e-18 M=1
c303 vdd n272 77.6e-18 M=1
c304 vdd n270 21.34e-18 M=1
c305 vdd n269 21.34e-18 M=1
c306 vdd n264 73.72e-18 M=1
c307 vdd n257 27.16e-18 M=1
c308 vdd n251 23.28e-18 M=1
c309 vdd n250 27.16e-18 M=1
c310 vdd n249 23.28e-18 M=1
c311 vdd n246 73.72e-18 M=1
c312 vdd n244 23.28e-18 M=1
c313 vdd n242 27.16e-18 M=1
c314 vdd n241 23.28e-18 M=1
c315 vdd n238 21.34e-18 M=1
c316 vdd n236 21.34e-18 M=1
c317 vdd n235 27.16e-18 M=1
c318 vdd n220 23.28e-18 M=1
c319 vdd n217 50.44e-18 M=1
c320 vdd n215 89.24e-18 M=1
c321 vdd n213 77.6e-18 M=1
c322 vdd n209 89.24e-18 M=1
c323 vdd n204 89.24e-18 M=1
c324 vdd n202 89.24e-18 M=1
c325 vdd n201 50.44e-18 M=1
c326 vdd n198 77.6e-18 M=1
c327 vdd n190 23.28e-18 M=1
c328 vdd n182 27.16e-18 M=1
c329 vdd n181 21.34e-18 M=1
c330 vdd n179 21.34e-18 M=1
c331 vdd n176 23.28e-18 M=1
c332 vdd n175 27.16e-18 M=1
c333 vdd n174 23.28e-18 M=1
c334 vdd n172 73.72e-18 M=1
c335 vdd n168 23.28e-18 M=1
c336 vdd n167 27.16e-18 M=1
c337 vdd n166 23.28e-18 M=1
c338 vdd n160 27.16e-18 M=1
c339 vdd n154 73.72e-18 M=1
c340 vdd n148 21.34e-18 M=1
c341 vdd n147 21.34e-18 M=1
c342 vdd n142 73.72e-18 M=1
c343 vdd n135 77.6e-18 M=1
c344 vdd n128 89.24e-18 M=1
c345 vdd n125 89.24e-18 M=1
c346 vdd n121 73.72e-18 M=1
c347 vdd n116 77.6e-18 M=1
c348 vdd n114 21.34e-18 M=1
c349 vdd n113 21.34e-18 M=1
c350 vdd n108 73.72e-18 M=1
c351 vdd n101 27.16e-18 M=1
c352 vdd n95 23.28e-18 M=1
c353 vdd n94 27.16e-18 M=1
c354 vdd n93 23.28e-18 M=1
c355 vdd n90 73.72e-18 M=1
c356 vdd n88 23.28e-18 M=1
c357 vdd n86 27.16e-18 M=1
c358 vdd n85 23.28e-18 M=1
c359 vdd n82 21.34e-18 M=1
c360 vdd n80 21.34e-18 M=1
c361 vdd n79 27.16e-18 M=1
c362 vdd n64 23.28e-18 M=1
c363 vdd n61 50.44e-18 M=1
c364 vdd n59 89.24e-18 M=1
c365 vdd n57 77.6e-18 M=1
c366 vdd n53 89.24e-18 M=1
c367 vdd a9 54.32e-18 M=1
c368 vdd a8 77.6e-18 M=1
c369 vdd a7 54.32e-18 M=1
c370 vdd a6 77.6e-18 M=1
c371 vdd a5 54.32e-18 M=1
c372 vdd a4 77.6e-18 M=1
c373 vdd a3 54.32e-18 M=1
c374 vdd a2 77.6e-18 M=1
c375 vdd a1 54.32e-18 M=1
c376 vdd a0 77.6e-18 M=1
c377 vdd b15 77.6e-18 M=1
c378 vdd b14 54.32e-18 M=1
c379 vdd b13 77.6e-18 M=1
c380 vdd b12 54.32e-18 M=1
c381 vdd b11 77.6e-18 M=1
c382 vdd b10 54.32e-18 M=1
c383 vdd a15 54.32e-18 M=1
c384 vdd a14 77.6e-18 M=1
c385 vdd a13 54.32e-18 M=1
c386 vdd a12 77.6e-18 M=1
c387 vdd a11 54.32e-18 M=1
c388 vdd a10 77.6e-18 M=1
c389 vdd cin 89.24e-18 M=1
c390 vdd b9 77.6e-18 M=1
c391 vdd b8 54.32e-18 M=1
c392 vdd b7 77.6e-18 M=1
c393 vdd b6 54.32e-18 M=1
c394 vdd b5 77.6e-18 M=1
c395 vdd b4 54.32e-18 M=1
c396 vdd b3 77.6e-18 M=1
c397 vdd b2 54.32e-18 M=1
c398 vdd b1 77.6e-18 M=1
c399 vdd b0 54.32e-18 M=1
c400 n356 n358 84.08e-18 M=1
c401 n354 n361 84.08e-18 M=1
c402 n353 n357 84.08e-18 M=1
c403 n350 n354 84.08e-18 M=1
c404 n348 n358 84.08e-18 M=1
c405 n346 n357 84.08e-18 M=1
c406 n345 n354 84.08e-18 M=1
c407 n344 n346 84.08e-18 M=1
c408 n342 n346 84.08e-18 M=1
c409 n335 n342 84.08e-18 M=1
c410 n328 n349 84.08e-18 M=1
c411 n328 n343 84.08e-18 M=1
c412 n328 n337 84.08e-18 M=1
c413 n327 n342 84.08e-18 M=1
c414 n318 n342 84.08e-18 M=1
c415 n303 n310 84.08e-18 M=1
c416 n298 n317 84.08e-18 M=1
c417 n298 n311 84.08e-18 M=1
c418 n298 n304 84.08e-18 M=1
c419 n297 n310 84.08e-18 M=1
c420 n291 n312 84.08e-18 M=1
c421 n291 n305 84.08e-18 M=1
c422 n290 n310 84.08e-18 M=1
c423 n284 n306 84.08e-18 M=1
c424 n284 n299 84.08e-18 M=1
c425 n276 n281 84.08e-18 M=1
c426 n272 n353 84.08e-18 M=1
c427 n269 n277 84.08e-18 M=1
c428 n268 n272 84.08e-18 M=1
c429 n267 n281 84.08e-18 M=1
c430 n264 n285 84.08e-18 M=1
c431 n264 n278 84.08e-18 M=1
c432 n264 n270 84.08e-18 M=1
c433 n263 n277 84.08e-18 M=1
c434 n261 n272 84.08e-18 M=1
c435 n256 n277 84.08e-18 M=1
c436 n236 n246 84.08e-18 M=1
c437 n232 n255 84.08e-18 M=1
c438 n232 n247 84.08e-18 M=1
c439 n232 n238 84.08e-18 M=1
c440 n231 n246 84.08e-18 M=1
c441 n225 n246 84.08e-18 M=1
c442 n221 n291 84.08e-18 M=1
c443 n220 n232 84.08e-18 M=1
c444 n220 n230 84.08e-18 M=1
c445 n217 n221 84.08e-18 M=1
c446 n217 n220 84.08e-18 M=1
c447 n213 n229 84.08e-18 M=1
c448 n213 n224 84.08e-18 M=1
c449 n212 n213 84.08e-18 M=1
c450 n209 n226 84.08e-18 M=1
c451 n209 n218 84.08e-18 M=1
c452 n204 n346 84.08e-18 M=1
c453 n200 n202 84.08e-18 M=1
c454 n198 n206 84.08e-18 M=1
c455 n197 n201 84.08e-18 M=1
c456 n194 n198 84.08e-18 M=1
c457 n192 n202 84.08e-18 M=1
c458 n190 n201 84.08e-18 M=1
c459 n189 n198 84.08e-18 M=1
c460 n188 n190 84.08e-18 M=1
c461 n186 n190 84.08e-18 M=1
c462 n179 n186 84.08e-18 M=1
c463 n172 n193 84.08e-18 M=1
c464 n172 n187 84.08e-18 M=1
c465 n172 n181 84.08e-18 M=1
c466 n171 n186 84.08e-18 M=1
c467 n162 n186 84.08e-18 M=1
c468 n147 n154 84.08e-18 M=1
c469 n142 n161 84.08e-18 M=1
c470 n142 n155 84.08e-18 M=1
c471 n142 n148 84.08e-18 M=1
c472 n141 n154 84.08e-18 M=1
c473 n135 n156 84.08e-18 M=1
c474 n135 n149 84.08e-18 M=1
c475 n134 n154 84.08e-18 M=1
c476 n128 n150 84.08e-18 M=1
c477 n128 n143 84.08e-18 M=1
c478 n120 n125 84.08e-18 M=1
c479 n116 n197 84.08e-18 M=1
c480 n113 n121 84.08e-18 M=1
c481 n112 n116 84.08e-18 M=1
c482 n111 n125 84.08e-18 M=1
c483 n108 n129 84.08e-18 M=1
c484 n108 n122 84.08e-18 M=1
c485 n108 n114 84.08e-18 M=1
c486 n107 n121 84.08e-18 M=1
c487 n105 n116 84.08e-18 M=1
c488 n100 n121 84.08e-18 M=1
c489 n80 n90 84.08e-18 M=1
c490 n76 n99 84.08e-18 M=1
c491 n76 n91 84.08e-18 M=1
c492 n76 n82 84.08e-18 M=1
c493 n75 n90 84.08e-18 M=1
c494 n69 n90 84.08e-18 M=1
c495 n65 n135 84.08e-18 M=1
c496 n64 n215 84.08e-18 M=1
c497 n64 n76 84.08e-18 M=1
c498 n64 n74 84.08e-18 M=1
c499 n61 n65 84.08e-18 M=1
c500 n61 n64 84.08e-18 M=1
c501 n59 n190 84.08e-18 M=1
c502 n57 n73 84.08e-18 M=1
c503 n57 n68 84.08e-18 M=1
c504 n56 n57 84.08e-18 M=1
c505 n53 n70 84.08e-18 M=1
c506 n53 n62 84.08e-18 M=1
c507 s2 n298 84.08e-18 M=1
c508 s2 n286 84.08e-18 M=1
c509 s2 n281 84.08e-18 M=1
c510 s2 n279 84.08e-18 M=1
c511 a9 n116 84.08e-18 M=1
c512 s1 n328 84.08e-18 M=1
c513 s1 n313 84.08e-18 M=1
c514 s1 n307 84.08e-18 M=1
c515 s1 n291 84.08e-18 M=1
c516 a8 n53 84.08e-18 M=1
c517 s0 n358 84.08e-18 M=1
c518 s0 n340 84.08e-18 M=1
c519 s0 n333 84.08e-18 M=1
c520 a7 n57 84.08e-18 M=1
c521 a6 n125 84.08e-18 M=1
c522 a5 n135 84.08e-18 M=1
c523 a4 n202 84.08e-18 M=1
c524 a3 n213 84.08e-18 M=1
c525 a2 n281 84.08e-18 M=1
c526 a1 n291 84.08e-18 M=1
c527 a0 n358 84.08e-18 M=1
c528 b15 n354 84.08e-18 M=1
c529 b14 n284 84.08e-18 M=1
c530 b13 n272 84.08e-18 M=1
c531 b12 n209 84.08e-18 M=1
c532 b11 n198 84.08e-18 M=1
c533 b10 n128 84.08e-18 M=1
c534 gnd n361 130.96e-18 M=1
c535 gnd n358 473.08e-18 M=1
c536 gnd n357 79.8e-18 M=1
c537 gnd n356 34.72e-18 M=1
c538 gnd n354 344.56e-18 M=1
c539 gnd n353 130.96e-18 M=1
c540 gnd n350 34.72e-18 M=1
c541 gnd n349 127.76e-18 M=1
c542 gnd n348 123.04e-18 M=1
c543 gnd n346 396.48e-18 M=1
c544 gnd n345 123.04e-18 M=1
c545 gnd n344 34.72e-18 M=1
c546 gnd n343 99.44e-18 M=1
c547 gnd n342 228.24e-18 M=1
c548 gnd n340 123.04e-18 M=1
c549 gnd n338 93.2e-18 M=1
c550 gnd n337 42.64e-18 M=1
c551 gnd n335 42.64e-18 M=1
c552 gnd n333 34.72e-18 M=1
c553 gnd n332 34.72e-18 M=1
c554 gnd n331 93.2e-18 M=1
c555 gnd n330 34.72e-18 M=1
c556 gnd n328 228.24e-18 M=1
c557 gnd n327 99.44e-18 M=1
c558 gnd n324 34.72e-18 M=1
c559 gnd n323 93.2e-18 M=1
c560 gnd n322 34.72e-18 M=1
c561 gnd n321 34.72e-18 M=1
c562 gnd n318 127.76e-18 M=1
c563 gnd n317 127.76e-18 M=1
c564 gnd n316 93.2e-18 M=1
c565 gnd n315 123.04e-18 M=1
c566 gnd n313 123.04e-18 M=1
c567 gnd n312 123.04e-18 M=1
c568 gnd n311 99.44e-18 M=1
c569 gnd n310 250.48e-18 M=1
c570 gnd n307 34.72e-18 M=1
c571 gnd n306 123.04e-18 M=1
c572 gnd n305 34.72e-18 M=1
c573 gnd n304 42.64e-18 M=1
c574 gnd n303 42.64e-18 M=1
c575 gnd n299 34.72e-18 M=1
c576 gnd n298 250.48e-18 M=1
c577 gnd n297 99.44e-18 M=1
c578 gnd n296 34.72e-18 M=1
c579 gnd n291 344.56e-18 M=1
c580 gnd n290 127.76e-18 M=1
c581 gnd n289 123.04e-18 M=1
c582 gnd n286 123.04e-18 M=1
c583 gnd n285 127.76e-18 M=1
c584 gnd n284 344.56e-18 M=1
c585 gnd n281 344.56e-18 M=1
c586 gnd n279 34.72e-18 M=1
c587 gnd n278 99.44e-18 M=1
c588 gnd n277 250.48e-18 M=1
c589 gnd n276 34.72e-18 M=1
c590 gnd n272 344.56e-18 M=1
c591 gnd n270 42.64e-18 M=1
c592 gnd n269 42.64e-18 M=1
c593 gnd n268 34.72e-18 M=1
c594 gnd n267 123.04e-18 M=1
c595 gnd n266 34.72e-18 M=1
c596 gnd n264 250.48e-18 M=1
c597 gnd n263 99.44e-18 M=1
c598 gnd n261 123.04e-18 M=1
c599 gnd n260 123.04e-18 M=1
c600 gnd n258 123.04e-18 M=1
c601 gnd n257 93.2e-18 M=1
c602 gnd n256 127.76e-18 M=1
c603 gnd n255 127.76e-18 M=1
c604 gnd n252 34.72e-18 M=1
c605 gnd n251 34.72e-18 M=1
c606 gnd n250 93.2e-18 M=1
c607 gnd n249 34.72e-18 M=1
c608 gnd n247 99.44e-18 M=1
c609 gnd n246 228.24e-18 M=1
c610 gnd n244 34.72e-18 M=1
c611 gnd n242 93.2e-18 M=1
c612 gnd n241 34.72e-18 M=1
c613 gnd n240 34.72e-18 M=1
c614 gnd n238 42.64e-18 M=1
c615 gnd n236 42.64e-18 M=1
c616 gnd n235 93.2e-18 M=1
c617 gnd n234 123.04e-18 M=1
c618 gnd n232 228.24e-18 M=1
c619 gnd n231 99.44e-18 M=1
c620 gnd n230 34.72e-18 M=1
c621 gnd n229 123.04e-18 M=1
c622 gnd n226 123.04e-18 M=1
c623 gnd n225 127.76e-18 M=1
c624 gnd n224 34.72e-18 M=1
c625 gnd n221 130.96e-18 M=1
c626 gnd n220 396.48e-18 M=1
c627 gnd n218 34.72e-18 M=1
c628 gnd n217 79.8e-18 M=1
c629 gnd n215 34.72e-18 M=1
c630 gnd n213 344.56e-18 M=1
c631 gnd n212 130.96e-18 M=1
c632 gnd n209 473.08e-18 M=1
c633 gnd n206 130.96e-18 M=1
c634 gnd n204 34.72e-18 M=1
c635 gnd n202 473.08e-18 M=1
c636 gnd n201 79.8e-18 M=1
c637 gnd n200 34.72e-18 M=1
c638 gnd n198 344.56e-18 M=1
c639 gnd n197 130.96e-18 M=1
c640 gnd n194 34.72e-18 M=1
c641 gnd n193 127.76e-18 M=1
c642 gnd n192 123.04e-18 M=1
c643 gnd n190 396.48e-18 M=1
c644 gnd n189 123.04e-18 M=1
c645 gnd n188 34.72e-18 M=1
c646 gnd n187 99.44e-18 M=1
c647 gnd n186 228.24e-18 M=1
c648 gnd n184 123.04e-18 M=1
c649 gnd n182 93.2e-18 M=1
c650 gnd n181 42.64e-18 M=1
c651 gnd n179 42.64e-18 M=1
c652 gnd n177 34.72e-18 M=1
c653 gnd n176 34.72e-18 M=1
c654 gnd n175 93.2e-18 M=1
c655 gnd n174 34.72e-18 M=1
c656 gnd n172 228.24e-18 M=1
c657 gnd n171 99.44e-18 M=1
c658 gnd n168 34.72e-18 M=1
c659 gnd n167 93.2e-18 M=1
c660 gnd n166 34.72e-18 M=1
c661 gnd n165 34.72e-18 M=1
c662 gnd n162 127.76e-18 M=1
c663 gnd n161 127.76e-18 M=1
c664 gnd n160 93.2e-18 M=1
c665 gnd n159 123.04e-18 M=1
c666 gnd n157 123.04e-18 M=1
c667 gnd n156 123.04e-18 M=1
c668 gnd n155 99.44e-18 M=1
c669 gnd n154 250.48e-18 M=1
c670 gnd n151 34.72e-18 M=1
c671 gnd n150 123.04e-18 M=1
c672 gnd n149 34.72e-18 M=1
c673 gnd n148 42.64e-18 M=1
c674 gnd n147 42.64e-18 M=1
c675 gnd n143 34.72e-18 M=1
c676 gnd n142 250.48e-18 M=1
c677 gnd n141 99.44e-18 M=1
c678 gnd n140 34.72e-18 M=1
c679 gnd n135 344.56e-18 M=1
c680 gnd n134 127.76e-18 M=1
c681 gnd n133 123.04e-18 M=1
c682 gnd n130 123.04e-18 M=1
c683 gnd n129 127.76e-18 M=1
c684 gnd n128 344.56e-18 M=1
c685 gnd n125 344.56e-18 M=1
c686 gnd n123 34.72e-18 M=1
c687 gnd n122 99.44e-18 M=1
c688 gnd n121 250.48e-18 M=1
c689 gnd n120 34.72e-18 M=1
c690 gnd n116 344.56e-18 M=1
c691 gnd n114 42.64e-18 M=1
c692 gnd n113 42.64e-18 M=1
c693 gnd n112 34.72e-18 M=1
c694 gnd n111 123.04e-18 M=1
c695 gnd n110 34.72e-18 M=1
c696 gnd n108 250.48e-18 M=1
c697 gnd n107 99.44e-18 M=1
c698 gnd n105 123.04e-18 M=1
c699 gnd n104 123.04e-18 M=1
c700 gnd n102 123.04e-18 M=1
c701 gnd n101 93.2e-18 M=1
c702 gnd n100 127.76e-18 M=1
c703 gnd n99 127.76e-18 M=1
c704 gnd n96 34.72e-18 M=1
c705 gnd n95 34.72e-18 M=1
c706 gnd n94 93.2e-18 M=1
c707 gnd n93 34.72e-18 M=1
c708 gnd n91 99.44e-18 M=1
c709 gnd n90 228.24e-18 M=1
c710 gnd n88 34.72e-18 M=1
c711 gnd n86 93.2e-18 M=1
c712 gnd n85 34.72e-18 M=1
c713 gnd n84 34.72e-18 M=1
c714 gnd n82 42.64e-18 M=1
c715 gnd n80 42.64e-18 M=1
c716 gnd n79 93.2e-18 M=1
c717 gnd n78 123.04e-18 M=1
c718 gnd n76 228.24e-18 M=1
c719 gnd n75 99.44e-18 M=1
c720 gnd n74 34.72e-18 M=1
c721 gnd n73 123.04e-18 M=1
c722 gnd n70 123.04e-18 M=1
c723 gnd n69 127.76e-18 M=1
c724 gnd n68 34.72e-18 M=1
c725 gnd n65 130.96e-18 M=1
c726 gnd n64 396.48e-18 M=1
c727 gnd n62 34.72e-18 M=1
c728 gnd n61 79.8e-18 M=1
c729 gnd n59 34.72e-18 M=1
c730 gnd n57 344.56e-18 M=1
c731 gnd n56 130.96e-18 M=1
c732 gnd n53 473.08e-18 M=1
c733 gnd s2 344.56e-18 M=1
c734 gnd a9 128.52e-18 M=1
c735 gnd s1 344.56e-18 M=1
c736 gnd s0 344.56e-18 M=1
c737 gnd a7 128.52e-18 M=1
c738 gnd a5 128.52e-18 M=1
c739 gnd a3 128.52e-18 M=1
c740 gnd a1 128.52e-18 M=1
c741 gnd b14 128.52e-18 M=1
c742 gnd b12 128.52e-18 M=1
c743 gnd b10 128.52e-18 M=1
c744 a15 n354 84.08e-18 M=1
c745 a15 gnd 128.52e-18 M=1
c746 a14 n284 84.08e-18 M=1
c747 a13 n272 84.08e-18 M=1
c748 a13 gnd 128.52e-18 M=1
c749 a12 n209 84.08e-18 M=1
c750 a11 n198 84.08e-18 M=1
c751 a11 gnd 128.52e-18 M=1
c752 a10 n128 84.08e-18 M=1
c753 cin n220 84.08e-18 M=1
c754 cin s0 84.08e-18 M=1
c755 s15 n354 84.08e-18 M=1
c756 s15 n321 84.08e-18 M=1
c757 s15 n315 84.08e-18 M=1
c758 s15 n310 84.08e-18 M=1
c759 s15 gnd 344.56e-18 M=1
c760 s14 n296 84.08e-18 M=1
c761 s14 n289 84.08e-18 M=1
c762 s14 n284 84.08e-18 M=1
c763 s14 n277 84.08e-18 M=1
c764 s14 gnd 344.56e-18 M=1
c765 s13 n272 84.08e-18 M=1
c766 s13 n266 84.08e-18 M=1
c767 s13 n260 84.08e-18 M=1
c768 s13 n246 84.08e-18 M=1
c769 s13 gnd 344.56e-18 M=1
c770 s12 n240 84.08e-18 M=1
c771 s12 n234 84.08e-18 M=1
c772 s12 n209 84.08e-18 M=1
c773 s12 n204 84.08e-18 M=1
c774 s12 gnd 344.56e-18 M=1
c775 s11 n198 84.08e-18 M=1
c776 s11 n165 84.08e-18 M=1
c777 s11 n159 84.08e-18 M=1
c778 s11 n154 84.08e-18 M=1
c779 s11 gnd 344.56e-18 M=1
c780 s10 n140 84.08e-18 M=1
c781 s10 n133 84.08e-18 M=1
c782 s10 n128 84.08e-18 M=1
c783 s10 n121 84.08e-18 M=1
c784 s10 gnd 344.56e-18 M=1
c785 cout gnd 34.72e-18 M=1
c786 b9 n116 84.08e-18 M=1
c787 b8 n53 84.08e-18 M=1
c788 b8 gnd 128.52e-18 M=1
c789 b7 n57 84.08e-18 M=1
c790 b6 n125 84.08e-18 M=1
c791 b6 gnd 128.52e-18 M=1
c792 b5 n135 84.08e-18 M=1
c793 b4 n202 84.08e-18 M=1
c794 b4 gnd 128.52e-18 M=1
c795 s9 n116 84.08e-18 M=1
c796 s9 n110 84.08e-18 M=1
c797 s9 n104 84.08e-18 M=1
c798 s9 n90 84.08e-18 M=1
c799 s9 gnd 344.56e-18 M=1
c800 b3 n213 84.08e-18 M=1
c801 s8 n84 84.08e-18 M=1
c802 s8 n78 84.08e-18 M=1
c803 s8 n59 84.08e-18 M=1
c804 s8 n53 84.08e-18 M=1
c805 s8 gnd 344.56e-18 M=1
c806 b2 n281 84.08e-18 M=1
c807 b2 gnd 128.52e-18 M=1
c808 s7 n108 84.08e-18 M=1
c809 s7 n102 84.08e-18 M=1
c810 s7 n96 84.08e-18 M=1
c811 s7 n57 84.08e-18 M=1
c812 s7 gnd 344.56e-18 M=1
c813 b1 n291 84.08e-18 M=1
c814 s6 n142 84.08e-18 M=1
c815 s6 n130 84.08e-18 M=1
c816 s6 n125 84.08e-18 M=1
c817 s6 n123 84.08e-18 M=1
c818 s6 gnd 344.56e-18 M=1
c819 b0 n358 84.08e-18 M=1
c820 b0 gnd 128.52e-18 M=1
c821 s5 n172 84.08e-18 M=1
c822 s5 n157 84.08e-18 M=1
c823 s5 n151 84.08e-18 M=1
c824 s5 n135 84.08e-18 M=1
c825 s5 gnd 344.56e-18 M=1
c826 vdd n435 29.32e-18 M=1
c827 vdd n434 58.64e-18 M=1
c828 vdd n433 58.64e-18 M=1
c829 vdd n432 58.64e-18 M=1
c830 vdd n431 58.64e-18 M=1
c831 vdd n430 58.64e-18 M=1
c832 vdd n429 58.64e-18 M=1
c833 vdd n428 29.32e-18 M=1
c834 vdd n427 29.32e-18 M=1
c835 vdd n426 58.64e-18 M=1
c836 vdd n425 58.64e-18 M=1
c837 vdd n424 58.64e-18 M=1
c838 vdd n423 58.64e-18 M=1
c839 vdd n422 58.64e-18 M=1
c840 vdd n421 58.64e-18 M=1
c841 vdd n420 29.32e-18 M=1
c842 vdd n361 69.44e-18 M=1
c843 vdd n358 53e-18 M=1
c844 vdd n357 60.76e-18 M=1
c845 vdd n356 34.72e-18 M=1
c846 vdd n354 34.72e-18 M=1
c847 vdd n353 69.44e-18 M=1
c848 vdd n350 34.72e-18 M=1
c849 vdd n349 34.72e-18 M=1
c850 vdd n348 56.96e-18 M=1
c851 vdd n346 34.72e-18 M=1
c852 vdd n345 56.96e-18 M=1
c853 vdd n344 34.72e-18 M=1
c854 vdd n343 34.72e-18 M=1
c855 vdd n342 69.44e-18 M=1
c856 vdd n340 56.96e-18 M=1
c857 vdd n338 61.68e-18 M=1
c858 vdd n337 42.64e-18 M=1
c859 vdd n335 42.64e-18 M=1
c860 vdd n333 34.72e-18 M=1
c861 vdd n332 34.72e-18 M=1
c862 vdd n331 61.68e-18 M=1
c863 vdd n330 34.72e-18 M=1
c864 vdd n328 69.44e-18 M=1
c865 vdd n327 34.72e-18 M=1
c866 vdd n324 34.72e-18 M=1
c867 vdd n323 61.68e-18 M=1
c868 vdd n322 34.72e-18 M=1
c869 vdd n321 34.72e-18 M=1
c870 vdd n318 34.72e-18 M=1
c871 vdd n317 34.72e-18 M=1
c872 vdd n316 61.68e-18 M=1
c873 vdd n315 56.96e-18 M=1
c874 vdd n313 56.96e-18 M=1
c875 vdd n312 56.96e-18 M=1
c876 vdd n311 34.72e-18 M=1
c877 vdd n310 124.72e-18 M=1
c878 vdd n307 34.72e-18 M=1
c879 vdd n306 56.96e-18 M=1
c880 vdd n305 34.72e-18 M=1
c881 vdd n304 42.64e-18 M=1
c882 vdd n303 42.64e-18 M=1
c883 vdd n299 34.72e-18 M=1
c884 vdd n298 124.72e-18 M=1
c885 vdd n297 34.72e-18 M=1
c886 vdd n296 34.72e-18 M=1
c887 vdd n291 34.72e-18 M=1
c888 vdd n290 34.72e-18 M=1
c889 vdd n289 56.96e-18 M=1
c890 vdd n286 56.96e-18 M=1
c891 vdd n285 34.72e-18 M=1
c892 vdd n284 34.72e-18 M=1
c893 vdd n281 34.72e-18 M=1
c894 vdd n279 34.72e-18 M=1
c895 vdd n278 34.72e-18 M=1
c896 vdd n277 124.72e-18 M=1
c897 vdd n276 34.72e-18 M=1
c898 vdd n272 34.72e-18 M=1
c899 vdd n270 42.64e-18 M=1
c900 vdd n269 42.64e-18 M=1
c901 vdd n268 34.72e-18 M=1
c902 vdd n267 56.96e-18 M=1
c903 vdd n266 34.72e-18 M=1
c904 vdd n264 124.72e-18 M=1
c905 vdd n263 34.72e-18 M=1
c906 vdd n261 56.96e-18 M=1
c907 vdd n260 56.96e-18 M=1
c908 vdd n258 56.96e-18 M=1
c909 vdd n257 61.68e-18 M=1
c910 vdd n256 34.72e-18 M=1
c911 vdd n255 34.72e-18 M=1
c912 vdd n252 34.72e-18 M=1
c913 vdd n251 34.72e-18 M=1
c914 vdd n250 61.68e-18 M=1
c915 vdd n249 34.72e-18 M=1
c916 vdd n247 34.72e-18 M=1
c917 vdd n246 69.44e-18 M=1
c918 vdd n244 34.72e-18 M=1
c919 vdd n242 61.68e-18 M=1
c920 vdd n241 34.72e-18 M=1
c921 vdd n240 34.72e-18 M=1
c922 vdd n238 42.64e-18 M=1
c923 vdd n236 42.64e-18 M=1
c924 vdd n235 61.68e-18 M=1
c925 vdd n234 56.96e-18 M=1
c926 vdd n232 69.44e-18 M=1
c927 vdd n231 34.72e-18 M=1
c928 vdd n230 34.72e-18 M=1
c929 vdd n229 56.96e-18 M=1
c930 vdd n226 56.96e-18 M=1
c931 vdd n225 34.72e-18 M=1
c932 vdd n224 34.72e-18 M=1
c933 vdd n221 69.44e-18 M=1
c934 vdd n220 34.72e-18 M=1
c935 vdd n218 34.72e-18 M=1
c936 vdd n217 60.76e-18 M=1
c937 vdd n215 34.72e-18 M=1
c938 vdd n213 34.72e-18 M=1
c939 vdd n212 69.44e-18 M=1
c940 vdd n209 53e-18 M=1
c941 vdd n206 69.44e-18 M=1
c942 vdd n204 34.72e-18 M=1
c943 vdd n202 53e-18 M=1
c944 vdd n201 60.76e-18 M=1
c945 vdd n200 34.72e-18 M=1
c946 vdd n198 34.72e-18 M=1
c947 vdd n197 69.44e-18 M=1
c948 vdd n194 34.72e-18 M=1
c949 vdd n193 34.72e-18 M=1
c950 vdd n192 56.96e-18 M=1
c951 vdd n190 34.72e-18 M=1
c952 vdd n189 56.96e-18 M=1
c953 vdd n188 34.72e-18 M=1
c954 vdd n187 34.72e-18 M=1
c955 vdd n186 69.44e-18 M=1
c956 vdd n184 56.96e-18 M=1
c957 vdd n182 61.68e-18 M=1
c958 vdd n181 42.64e-18 M=1
c959 vdd n179 42.64e-18 M=1
c960 vdd n177 34.72e-18 M=1
c961 vdd n176 34.72e-18 M=1
c962 vdd n175 61.68e-18 M=1
c963 vdd n174 34.72e-18 M=1
c964 vdd n172 69.44e-18 M=1
c965 vdd n171 34.72e-18 M=1
c966 vdd n168 34.72e-18 M=1
c967 vdd n167 61.68e-18 M=1
c968 vdd n166 34.72e-18 M=1
c969 vdd n165 34.72e-18 M=1
c970 vdd n162 34.72e-18 M=1
c971 vdd n161 34.72e-18 M=1
c972 vdd n160 61.68e-18 M=1
c973 vdd n159 56.96e-18 M=1
c974 vdd n157 56.96e-18 M=1
c975 vdd n156 56.96e-18 M=1
c976 vdd n155 34.72e-18 M=1
c977 vdd n154 124.72e-18 M=1
c978 vdd n151 34.72e-18 M=1
c979 vdd n150 56.96e-18 M=1
c980 vdd n149 34.72e-18 M=1
c981 vdd n148 42.64e-18 M=1
c982 vdd n147 42.64e-18 M=1
c983 vdd n143 34.72e-18 M=1
c984 vdd n142 124.72e-18 M=1
c985 vdd n141 34.72e-18 M=1
c986 vdd n140 34.72e-18 M=1
c987 vdd n135 34.72e-18 M=1
c988 vdd n134 34.72e-18 M=1
c989 vdd n133 56.96e-18 M=1
c990 vdd n130 56.96e-18 M=1
c991 vdd n129 34.72e-18 M=1
c992 vdd n128 34.72e-18 M=1
c993 vdd n125 34.72e-18 M=1
c994 vdd n123 34.72e-18 M=1
c995 vdd n122 34.72e-18 M=1
c996 vdd n121 124.72e-18 M=1
c997 vdd n120 34.72e-18 M=1
c998 vdd n116 34.72e-18 M=1
c999 vdd n114 42.64e-18 M=1
c1000 vdd n113 42.64e-18 M=1
c1001 vdd n112 34.72e-18 M=1
c1002 vdd n111 56.96e-18 M=1
c1003 vdd n110 34.72e-18 M=1
c1004 vdd n108 124.72e-18 M=1
c1005 vdd n107 34.72e-18 M=1
c1006 vdd n105 56.96e-18 M=1
c1007 vdd n104 56.96e-18 M=1
c1008 vdd n102 56.96e-18 M=1
c1009 vdd n101 61.68e-18 M=1
c1010 vdd n100 34.72e-18 M=1
c1011 vdd n99 34.72e-18 M=1
c1012 vdd n96 34.72e-18 M=1
c1013 vdd n95 34.72e-18 M=1
c1014 vdd n94 61.68e-18 M=1
c1015 vdd n93 34.72e-18 M=1
c1016 vdd n91 34.72e-18 M=1
c1017 vdd n90 69.44e-18 M=1
c1018 vdd n88 34.72e-18 M=1
c1019 vdd n86 61.68e-18 M=1
c1020 vdd n85 34.72e-18 M=1
c1021 vdd n84 34.72e-18 M=1
c1022 vdd n82 42.64e-18 M=1
c1023 vdd n80 42.64e-18 M=1
c1024 vdd n79 61.68e-18 M=1
c1025 vdd n78 56.96e-18 M=1
c1026 vdd n76 69.44e-18 M=1
c1027 vdd n75 34.72e-18 M=1
c1028 vdd n74 34.72e-18 M=1
c1029 vdd n73 56.96e-18 M=1
c1030 vdd n70 56.96e-18 M=1
c1031 vdd n69 34.72e-18 M=1
c1032 vdd n68 34.72e-18 M=1
c1033 vdd n65 69.44e-18 M=1
c1034 vdd n64 34.72e-18 M=1
c1035 vdd n62 34.72e-18 M=1
c1036 vdd n61 60.76e-18 M=1
c1037 vdd n59 34.72e-18 M=1
c1038 vdd n57 34.72e-18 M=1
c1039 vdd n56 69.44e-18 M=1
c1040 vdd n53 53e-18 M=1
c1041 vdd s2 34.72e-18 M=1
c1042 vdd s1 34.72e-18 M=1
c1043 vdd s0 34.72e-18 M=1
c1044 vdd gnd 11.088e-15 M=1
c1045 vdd s15 34.72e-18 M=1
c1046 vdd s14 34.72e-18 M=1
c1047 vdd s13 34.72e-18 M=1
c1048 vdd s12 34.72e-18 M=1
c1049 vdd s11 34.72e-18 M=1
c1050 vdd s10 34.72e-18 M=1
c1051 vdd cout 34.72e-18 M=1
c1052 vdd s9 34.72e-18 M=1
c1053 vdd s8 34.72e-18 M=1
c1054 vdd s7 34.72e-18 M=1
c1055 vdd s6 34.72e-18 M=1
c1056 vdd s5 34.72e-18 M=1
c1057 s4 n215 84.08e-18 M=1
c1058 s4 n202 84.08e-18 M=1
c1059 s4 n184 84.08e-18 M=1
c1060 s4 n177 84.08e-18 M=1
c1061 s4 gnd 344.56e-18 M=1
c1062 s4 vdd 34.72e-18 M=1
c1063 s3 n264 84.08e-18 M=1
c1064 s3 n258 84.08e-18 M=1
c1065 s3 n252 84.08e-18 M=1
c1066 s3 n213 84.08e-18 M=1
c1067 s3 gnd 344.56e-18 M=1
c1068 s3 vdd 34.72e-18 M=1
c1069 n358 n419 85.36e-18 M=1
c1070 n358 n412 46.88e-18 M=1
c1071 n357 n416 46.88e-18 M=1
c1072 n356 n419 46.88e-18 M=1
c1073 n356 n358 83.84e-18 M=1
c1074 n354 n417 85.36e-18 M=1
c1075 n354 n413 46.88e-18 M=1
c1076 n350 n417 46.88e-18 M=1
c1077 n350 n354 83.84e-18 M=1
c1078 n348 n419 46.88e-18 M=1
c1079 n348 n358 83.84e-18 M=1
c1080 n348 n356 46.88e-18 M=1
c1081 n346 n416 85.36e-18 M=1
c1082 n346 n357 83.84e-18 M=1
c1083 n345 n417 46.88e-18 M=1
c1084 n345 n354 83.84e-18 M=1
c1085 n345 n350 46.88e-18 M=1
c1086 n344 n416 46.88e-18 M=1
c1087 n344 n357 178.17e-18 M=1
c1088 n344 n346 83.84e-18 M=1
c1089 n343 n349 46.88e-18 M=1
c1090 n342 n416 46.88e-18 M=1
c1091 n342 n357 93.76e-18 M=1
c1092 n342 n346 83.84e-18 M=1
c1093 n342 n344 46.88e-18 M=1
c1094 n340 n412 46.88e-18 M=1
c1095 n340 n358 46.88e-18 M=1
c1096 n339 n342 85.36e-18 M=1
c1097 n337 n349 46.88e-18 M=1
c1098 n337 n343 46.88e-18 M=1
c1099 n335 n342 83.84e-18 M=1
c1100 n335 n339 46.88e-18 M=1
c1101 n333 n412 46.88e-18 M=1
c1102 n333 n358 46.88e-18 M=1
c1103 n333 n340 46.88e-18 M=1
c1104 n328 n408 46.88e-18 M=1
c1105 n328 n343 83.84e-18 M=1
c1106 n328 n337 83.84e-18 M=1
c1107 n328 n330 46.88e-18 M=1
c1108 n327 n342 83.84e-18 M=1
c1109 n327 n335 46.88e-18 M=1
c1110 n325 n349 46.88e-18 M=1
c1111 n325 n337 46.88e-18 M=1
c1112 n325 n328 85.36e-18 M=1
c1113 n321 n413 46.88e-18 M=1
c1114 n321 n354 46.88e-18 M=1
c1115 n318 n339 46.88e-18 M=1
c1116 n318 n335 46.88e-18 M=1
c1117 n318 n327 46.88e-18 M=1
c1118 n317 n328 84.41e-18 M=1
c1119 n315 n413 46.88e-18 M=1
c1120 n315 n354 46.88e-18 M=1
c1121 n315 n321 46.88e-18 M=1
c1122 n313 n408 46.88e-18 M=1
c1123 n313 n328 46.88e-18 M=1
c1124 n312 n407 46.88e-18 M=1
c1125 n311 n328 84.41e-18 M=1
c1126 n311 n317 46.88e-18 M=1
c1127 n310 n413 46.88e-18 M=1
c1128 n310 n354 177.6e-18 M=1
c1129 n310 n327 84.41e-18 M=1
c1130 n310 n324 46.88e-18 M=1
c1131 n310 n321 131.29e-18 M=1
c1132 n310 n318 84.41e-18 M=1
c1133 n310 n315 46.88e-18 M=1
c1134 n309 n310 85.36e-18 M=1
c1135 n307 n408 46.88e-18 M=1
c1136 n307 n328 131.29e-18 M=1
c1137 n307 n313 46.88e-18 M=1
c1138 n306 n406 46.88e-18 M=1
c1139 n305 n407 46.88e-18 M=1
c1140 n305 n312 46.88e-18 M=1
c1141 n304 n317 46.88e-18 M=1
c1142 n304 n311 46.88e-18 M=1
c1143 n303 n310 83.84e-18 M=1
c1144 n303 n309 46.88e-18 M=1
c1145 n299 n406 46.88e-18 M=1
c1146 n299 n306 46.88e-18 M=1
c1147 n298 n401 46.88e-18 M=1
c1148 n298 n311 83.84e-18 M=1
c1149 n298 n304 83.84e-18 M=1
c1150 n297 n310 83.84e-18 M=1
c1151 n297 n303 46.88e-18 M=1
c1152 n296 n410 46.88e-18 M=1
c1153 n294 n317 46.88e-18 M=1
c1154 n294 n304 46.88e-18 M=1
c1155 n294 n298 85.36e-18 M=1
c1156 n291 n408 46.88e-18 M=1
c1157 n291 n407 85.36e-18 M=1
c1158 n291 n328 93.76e-18 M=1
c1159 n291 n317 83.84e-18 M=1
c1160 n291 n313 46.88e-18 M=1
c1161 n291 n312 83.84e-18 M=1
c1162 n291 n307 46.88e-18 M=1
c1163 n291 n305 83.84e-18 M=1
c1164 n290 n309 46.88e-18 M=1
c1165 n290 n303 46.88e-18 M=1
c1166 n290 n297 46.88e-18 M=1
c1167 n289 n410 46.88e-18 M=1
c1168 n289 n296 46.88e-18 M=1
c1169 n286 n401 46.88e-18 M=1
c1170 n286 n298 46.88e-18 M=1
c1171 n285 n298 84.41e-18 M=1
c1172 n284 n410 46.88e-18 M=1
c1173 n284 n406 85.36e-18 M=1
c1174 n284 n306 83.84e-18 M=1
c1175 n284 n299 83.84e-18 M=1
c1176 n284 n296 46.88e-18 M=1
c1177 n284 n289 46.88e-18 M=1
c1178 n281 n405 85.36e-18 M=1
c1179 n281 n401 46.88e-18 M=1
c1180 n281 n298 93.76e-18 M=1
c1181 n281 n286 46.88e-18 M=1
c1182 n279 n401 46.88e-18 M=1
c1183 n279 n298 131.29e-18 M=1
c1184 n279 n286 46.88e-18 M=1
c1185 n279 n281 46.88e-18 M=1
c1186 n278 n298 84.41e-18 M=1
c1187 n278 n285 46.88e-18 M=1
c1188 n277 n410 46.88e-18 M=1
c1189 n277 n322 46.88e-18 M=1
c1190 n277 n297 84.41e-18 M=1
c1191 n277 n296 131.29e-18 M=1
c1192 n277 n290 84.41e-18 M=1
c1193 n277 n289 46.88e-18 M=1
c1194 n277 n284 93.76e-18 M=1
c1195 n276 n405 46.88e-18 M=1
c1196 n276 n281 83.84e-18 M=1
c1197 n274 n277 85.36e-18 M=1
c1198 n272 n403 85.36e-18 M=1
c1199 n272 n402 46.88e-18 M=1
c1200 n270 n285 46.88e-18 M=1
c1201 n270 n278 46.88e-18 M=1
c1202 n269 n277 83.84e-18 M=1
c1203 n269 n274 46.88e-18 M=1
c1204 n268 n403 46.88e-18 M=1
c1205 n268 n272 83.84e-18 M=1
c1206 n267 n405 46.88e-18 M=1
c1207 n267 n281 83.84e-18 M=1
c1208 n267 n276 46.88e-18 M=1
c1209 n266 n402 46.88e-18 M=1
c1210 n266 n272 46.88e-18 M=1
c1211 n264 n397 46.88e-18 M=1
c1212 n264 n278 83.84e-18 M=1
c1213 n264 n270 83.84e-18 M=1
c1214 n263 n277 83.84e-18 M=1
c1215 n263 n269 46.88e-18 M=1
c1216 n262 n285 46.88e-18 M=1
c1217 n262 n270 46.88e-18 M=1
c1218 n262 n264 85.36e-18 M=1
c1219 n261 n403 46.88e-18 M=1
c1220 n261 n272 83.84e-18 M=1
c1221 n261 n268 46.88e-18 M=1
c1222 n260 n402 46.88e-18 M=1
c1223 n260 n272 46.88e-18 M=1
c1224 n260 n266 46.88e-18 M=1
c1225 n258 n397 46.88e-18 M=1
c1226 n258 n264 46.88e-18 M=1
c1227 n256 n274 46.88e-18 M=1
c1228 n256 n272 83.84e-18 M=1
c1229 n256 n269 46.88e-18 M=1
c1230 n256 n263 46.88e-18 M=1
c1231 n255 n264 84.41e-18 M=1
c1232 n252 n397 46.88e-18 M=1
c1233 n252 n264 131.29e-18 M=1
c1234 n252 n258 46.88e-18 M=1
c1235 n251 n298 46.88e-18 M=1
c1236 n249 n264 46.88e-18 M=1
c1237 n247 n264 84.41e-18 M=1
c1238 n247 n255 46.88e-18 M=1
c1239 n246 n402 46.88e-18 M=1
c1240 n246 n272 93.76e-18 M=1
c1241 n246 n266 131.29e-18 M=1
c1242 n246 n263 84.41e-18 M=1
c1243 n246 n260 46.88e-18 M=1
c1244 n246 n256 84.41e-18 M=1
c1245 n244 n246 46.88e-18 M=1
c1246 n243 n246 85.36e-18 M=1
c1247 n240 n398 46.88e-18 M=1
c1248 n238 n255 46.88e-18 M=1
c1249 n238 n247 46.88e-18 M=1
c1250 n236 n246 83.84e-18 M=1
c1251 n236 n243 46.88e-18 M=1
c1252 n234 n398 46.88e-18 M=1
c1253 n234 n240 46.88e-18 M=1
c1254 n232 n395 46.88e-18 M=1
c1255 n232 n247 83.84e-18 M=1
c1256 n232 n238 83.84e-18 M=1
c1257 n231 n246 83.84e-18 M=1
c1258 n231 n236 46.88e-18 M=1
c1259 n230 n395 46.88e-18 M=1
c1260 n230 n232 46.88e-18 M=1
c1261 n229 n393 46.88e-18 M=1
c1262 n228 n255 46.88e-18 M=1
c1263 n228 n238 46.88e-18 M=1
c1264 n228 n232 85.36e-18 M=1
c1265 n226 n392 46.88e-18 M=1
c1266 n225 n243 46.88e-18 M=1
c1267 n225 n236 46.88e-18 M=1
c1268 n225 n231 46.88e-18 M=1
c1269 n224 n393 46.88e-18 M=1
c1270 n224 n229 46.88e-18 M=1
c1271 n220 n395 85.36e-18 M=1
c1272 n220 n232 83.84e-18 M=1
c1273 n220 n230 83.84e-18 M=1
c1274 n218 n392 46.88e-18 M=1
c1275 n218 n226 46.88e-18 M=1
c1276 n217 n395 46.88e-18 M=1
c1277 n217 n232 93.76e-18 M=1
c1278 n217 n230 178.17e-18 M=1
c1279 n217 n220 83.84e-18 M=1
c1280 n215 n384 46.88e-18 M=1
c1281 n215 n367 46.88e-18 M=1
c1282 n213 n397 46.88e-18 M=1
c1283 n213 n393 85.36e-18 M=1
c1284 n213 n264 177.6e-18 M=1
c1285 n213 n258 46.88e-18 M=1
c1286 n213 n252 46.88e-18 M=1
c1287 n213 n229 83.84e-18 M=1
c1288 n213 n224 83.84e-18 M=1
c1289 n209 n398 46.88e-18 M=1
c1290 n209 n392 85.36e-18 M=1
c1291 n209 n240 46.88e-18 M=1
c1292 n209 n234 46.88e-18 M=1
c1293 n209 n226 83.84e-18 M=1
c1294 n209 n218 83.84e-18 M=1
c1295 n204 n416 46.88e-18 M=1
c1296 n204 n398 46.88e-18 M=1
c1297 n204 n357 46.88e-18 M=1
c1298 n204 n344 46.88e-18 M=1
c1299 n204 n342 46.88e-18 M=1
c1300 n204 n241 46.88e-18 M=1
c1301 n204 n240 131.29e-18 M=1
c1302 n204 n234 46.88e-18 M=1
c1303 n204 n231 84.6e-18 M=1
c1304 n204 n225 84.6e-18 M=1
c1305 n204 n209 93.76e-18 M=1
c1306 n202 n391 85.36e-18 M=1
c1307 n202 n384 46.88e-18 M=1
c1308 n202 n215 93.76e-18 M=1
c1309 n201 n388 46.88e-18 M=1
c1310 n200 n391 46.88e-18 M=1
c1311 n200 n202 83.84e-18 M=1
c1312 n198 n389 85.36e-18 M=1
c1313 n198 n385 46.88e-18 M=1
c1314 n194 n389 46.88e-18 M=1
c1315 n194 n198 83.84e-18 M=1
c1316 n193 n215 84.6e-18 M=1
c1317 n192 n391 46.88e-18 M=1
c1318 n192 n202 83.84e-18 M=1
c1319 n192 n200 46.88e-18 M=1
c1320 n190 n388 85.36e-18 M=1
c1321 n190 n201 83.84e-18 M=1
c1322 n189 n389 46.88e-18 M=1
c1323 n189 n198 83.84e-18 M=1
c1324 n189 n194 46.88e-18 M=1
c1325 n188 n388 46.88e-18 M=1
c1326 n188 n201 178.17e-18 M=1
c1327 n188 n190 83.84e-18 M=1
c1328 n187 n215 84.6e-18 M=1
c1329 n187 n193 46.88e-18 M=1
c1330 n186 n388 46.88e-18 M=1
c1331 n186 n201 93.76e-18 M=1
c1332 n186 n190 83.84e-18 M=1
c1333 n186 n188 46.88e-18 M=1
c1334 n184 n384 46.88e-18 M=1
c1335 n184 n215 46.88e-18 M=1
c1336 n184 n202 46.88e-18 M=1
c1337 n183 n186 85.36e-18 M=1
c1338 n181 n193 46.88e-18 M=1
c1339 n181 n187 46.88e-18 M=1
c1340 n179 n186 83.84e-18 M=1
c1341 n179 n183 46.88e-18 M=1
c1342 n177 n384 46.88e-18 M=1
c1343 n177 n215 131.29e-18 M=1
c1344 n177 n202 46.88e-18 M=1
c1345 n177 n184 46.88e-18 M=1
c1346 n176 n215 46.88e-18 M=1
c1347 n172 n380 46.88e-18 M=1
c1348 n172 n187 83.84e-18 M=1
c1349 n172 n181 83.84e-18 M=1
c1350 n172 n174 46.88e-18 M=1
c1351 n171 n186 83.84e-18 M=1
c1352 n171 n179 46.88e-18 M=1
c1353 n169 n193 46.88e-18 M=1
c1354 n169 n181 46.88e-18 M=1
c1355 n169 n172 85.36e-18 M=1
c1356 n165 n385 46.88e-18 M=1
c1357 n165 n198 46.88e-18 M=1
c1358 n162 n183 46.88e-18 M=1
c1359 n162 n179 46.88e-18 M=1
c1360 n162 n171 46.88e-18 M=1
c1361 n161 n172 84.41e-18 M=1
c1362 n159 n385 46.88e-18 M=1
c1363 n159 n198 46.88e-18 M=1
c1364 n159 n165 46.88e-18 M=1
c1365 n157 n380 46.88e-18 M=1
c1366 n157 n172 46.88e-18 M=1
c1367 n156 n379 46.88e-18 M=1
c1368 n155 n172 84.41e-18 M=1
c1369 n155 n161 46.88e-18 M=1
c1370 n154 n385 46.88e-18 M=1
c1371 n154 n198 177.6e-18 M=1
c1372 n154 n171 84.41e-18 M=1
c1373 n154 n168 46.88e-18 M=1
c1374 n154 n165 131.29e-18 M=1
c1375 n154 n162 84.41e-18 M=1
c1376 n154 n159 46.88e-18 M=1
c1377 n153 n154 85.36e-18 M=1
c1378 n151 n380 46.88e-18 M=1
c1379 n151 n172 131.29e-18 M=1
c1380 n151 n157 46.88e-18 M=1
c1381 n150 n378 46.88e-18 M=1
c1382 n149 n379 46.88e-18 M=1
c1383 n149 n156 46.88e-18 M=1
c1384 n148 n161 46.88e-18 M=1
c1385 n148 n155 46.88e-18 M=1
c1386 n147 n154 83.84e-18 M=1
c1387 n147 n153 46.88e-18 M=1
c1388 n143 n378 46.88e-18 M=1
c1389 n143 n150 46.88e-18 M=1
c1390 n142 n373 46.88e-18 M=1
c1391 n142 n155 83.84e-18 M=1
c1392 n142 n148 83.84e-18 M=1
c1393 n141 n154 83.84e-18 M=1
c1394 n141 n147 46.88e-18 M=1
c1395 n140 n382 46.88e-18 M=1
c1396 n138 n161 46.88e-18 M=1
c1397 n138 n148 46.88e-18 M=1
c1398 n138 n142 85.36e-18 M=1
c1399 n135 n380 46.88e-18 M=1
c1400 n135 n379 85.36e-18 M=1
c1401 n135 n172 93.76e-18 M=1
c1402 n135 n161 83.84e-18 M=1
c1403 n135 n157 46.88e-18 M=1
c1404 n135 n156 83.84e-18 M=1
c1405 n135 n151 46.88e-18 M=1
c1406 n135 n149 83.84e-18 M=1
c1407 n134 n153 46.88e-18 M=1
c1408 n134 n147 46.88e-18 M=1
c1409 n134 n141 46.88e-18 M=1
c1410 n133 n382 46.88e-18 M=1
c1411 n133 n140 46.88e-18 M=1
c1412 n130 n373 46.88e-18 M=1
c1413 n130 n142 46.88e-18 M=1
c1414 n129 n142 84.41e-18 M=1
c1415 n128 n382 46.88e-18 M=1
c1416 n128 n378 85.36e-18 M=1
c1417 n128 n150 83.84e-18 M=1
c1418 n128 n143 83.84e-18 M=1
c1419 n128 n140 46.88e-18 M=1
c1420 n128 n133 46.88e-18 M=1
c1421 n125 n377 85.36e-18 M=1
c1422 n125 n373 46.88e-18 M=1
c1423 n125 n142 93.76e-18 M=1
c1424 n125 n130 46.88e-18 M=1
c1425 n123 n373 46.88e-18 M=1
c1426 n123 n142 131.29e-18 M=1
c1427 n123 n130 46.88e-18 M=1
c1428 n123 n125 46.88e-18 M=1
c1429 n122 n142 84.41e-18 M=1
c1430 n122 n129 46.88e-18 M=1
c1431 n121 n382 46.88e-18 M=1
c1432 n121 n166 46.88e-18 M=1
c1433 n121 n141 84.41e-18 M=1
c1434 n121 n140 131.29e-18 M=1
c1435 n121 n134 84.41e-18 M=1
c1436 n121 n133 46.88e-18 M=1
c1437 n121 n128 93.76e-18 M=1
c1438 n120 n377 46.88e-18 M=1
c1439 n120 n125 83.84e-18 M=1
c1440 n118 n121 85.36e-18 M=1
c1441 n116 n375 85.36e-18 M=1
c1442 n116 n374 46.88e-18 M=1
c1443 n114 n129 46.88e-18 M=1
c1444 n114 n122 46.88e-18 M=1
c1445 n113 n121 83.84e-18 M=1
c1446 n113 n118 46.88e-18 M=1
c1447 n112 n375 46.88e-18 M=1
c1448 n112 n116 83.84e-18 M=1
c1449 n111 n377 46.88e-18 M=1
c1450 n111 n125 83.84e-18 M=1
c1451 n111 n120 46.88e-18 M=1
c1452 n110 n374 46.88e-18 M=1
c1453 n110 n116 46.88e-18 M=1
c1454 n108 n369 46.88e-18 M=1
c1455 n108 n122 83.84e-18 M=1
c1456 n108 n114 83.84e-18 M=1
c1457 n107 n121 83.84e-18 M=1
c1458 n107 n113 46.88e-18 M=1
c1459 n106 n129 46.88e-18 M=1
c1460 n106 n114 46.88e-18 M=1
c1461 n106 n108 85.36e-18 M=1
c1462 n105 n375 46.88e-18 M=1
c1463 n105 n116 83.84e-18 M=1
c1464 n105 n112 46.88e-18 M=1
c1465 n104 n374 46.88e-18 M=1
c1466 n104 n116 46.88e-18 M=1
c1467 n104 n110 46.88e-18 M=1
c1468 n102 n369 46.88e-18 M=1
c1469 n102 n108 46.88e-18 M=1
c1470 n100 n118 46.88e-18 M=1
c1471 n100 n116 83.84e-18 M=1
c1472 n100 n113 46.88e-18 M=1
c1473 n100 n107 46.88e-18 M=1
c1474 n99 n108 84.41e-18 M=1
c1475 n96 n369 46.88e-18 M=1
c1476 n96 n108 131.29e-18 M=1
c1477 n96 n102 46.88e-18 M=1
c1478 n95 n142 46.88e-18 M=1
c1479 n93 n108 46.88e-18 M=1
c1480 n91 n108 84.41e-18 M=1
c1481 n91 n99 46.88e-18 M=1
c1482 n90 n374 46.88e-18 M=1
c1483 n90 n116 93.76e-18 M=1
c1484 n90 n110 131.29e-18 M=1
c1485 n90 n107 84.41e-18 M=1
c1486 n90 n104 46.88e-18 M=1
c1487 n90 n100 84.41e-18 M=1
c1488 n88 n90 46.88e-18 M=1
c1489 n87 n90 85.36e-18 M=1
c1490 n84 n370 46.88e-18 M=1
c1491 n82 n99 46.88e-18 M=1
c1492 n82 n91 46.88e-18 M=1
c1493 n80 n90 83.84e-18 M=1
c1494 n80 n87 46.88e-18 M=1
c1495 n78 n370 46.88e-18 M=1
c1496 n78 n84 46.88e-18 M=1
c1497 n76 n367 46.88e-18 M=1
c1498 n76 n215 46.88e-18 M=1
c1499 n76 n91 83.84e-18 M=1
c1500 n76 n82 83.84e-18 M=1
c1501 n75 n90 83.84e-18 M=1
c1502 n75 n80 46.88e-18 M=1
c1503 n74 n367 46.88e-18 M=1
c1504 n74 n215 46.88e-18 M=1
c1505 n74 n76 46.88e-18 M=1
c1506 n73 n365 46.88e-18 M=1
c1507 n72 n99 46.88e-18 M=1
c1508 n72 n82 46.88e-18 M=1
c1509 n72 n76 85.36e-18 M=1
c1510 n70 n364 46.88e-18 M=1
c1511 n69 n87 46.88e-18 M=1
c1512 n69 n80 46.88e-18 M=1
c1513 n69 n75 46.88e-18 M=1
c1514 n68 n365 46.88e-18 M=1
c1515 n68 n73 46.88e-18 M=1
c1516 n64 n367 85.36e-18 M=1
c1517 n64 n76 83.84e-18 M=1
c1518 n64 n74 83.84e-18 M=1
c1519 n62 n364 46.88e-18 M=1
c1520 n62 n70 46.88e-18 M=1
c1521 n61 n367 46.88e-18 M=1
c1522 n61 n215 46.88e-18 M=1
c1523 n61 n76 93.76e-18 M=1
c1524 n61 n74 178.17e-18 M=1
c1525 n61 n64 83.84e-18 M=1
c1526 n59 n388 46.88e-18 M=1
c1527 n59 n370 46.88e-18 M=1
c1528 n59 n201 46.88e-18 M=1
c1529 n59 n188 46.88e-18 M=1
c1530 n59 n186 46.88e-18 M=1
c1531 n59 n85 46.88e-18 M=1
c1532 n59 n84 131.29e-18 M=1
c1533 n59 n78 46.88e-18 M=1
c1534 n59 n75 84.6e-18 M=1
c1535 n59 n69 84.6e-18 M=1
c1536 n57 n369 46.88e-18 M=1
c1537 n57 n365 85.36e-18 M=1
c1538 n57 n108 177.6e-18 M=1
c1539 n57 n102 46.88e-18 M=1
c1540 n57 n96 46.88e-18 M=1
c1541 n57 n73 83.84e-18 M=1
c1542 n57 n68 83.84e-18 M=1
c1543 n53 n370 46.88e-18 M=1
c1544 n53 n364 85.36e-18 M=1
c1545 n53 n84 46.88e-18 M=1
c1546 n53 n78 46.88e-18 M=1
c1547 n53 n70 83.84e-18 M=1
c1548 n53 n62 83.84e-18 M=1
c1549 n53 n59 93.76e-18 M=1
c1550 s2 n401 85.36e-18 M=1
c1551 s2 n286 83.84e-18 M=1
c1552 s2 n281 83.84e-18 M=1
c1553 s2 n279 83.84e-18 M=1
c1554 a9 n375 46.88e-18 M=1
c1555 a9 n116 83.84e-18 M=1
c1556 a9 n112 46.88e-18 M=1
c1557 a9 n105 46.88e-18 M=1
c1558 a9 n94 46.88e-18 M=1
c1559 s1 n408 85.36e-18 M=1
c1560 s1 n313 83.84e-18 M=1
c1561 s1 n307 83.84e-18 M=1
c1562 s1 n291 83.84e-18 M=1
c1563 a8 n364 46.88e-18 M=1
c1564 a8 n70 131.29e-18 M=1
c1565 a8 n62 131.29e-18 M=1
c1566 s0 n412 85.36e-18 M=1
c1567 s0 n358 83.84e-18 M=1
c1568 s0 n340 83.84e-18 M=1
c1569 s0 n333 83.84e-18 M=1
c1570 a7 n365 46.88e-18 M=1
c1571 a7 n86 46.88e-18 M=1
c1572 a7 n73 46.88e-18 M=1
c1573 a7 n68 46.88e-18 M=1
c1574 a7 n57 83.84e-18 M=1
c1575 a6 n377 46.88e-18 M=1
c1576 a6 n120 131.29e-18 M=1
c1577 a6 n111 131.29e-18 M=1
c1578 a5 n379 46.88e-18 M=1
c1579 a5 n167 46.88e-18 M=1
c1580 a5 n156 46.88e-18 M=1
c1581 a5 n149 46.88e-18 M=1
c1582 a5 n135 83.84e-18 M=1
c1583 a4 n391 46.88e-18 M=1
c1584 a4 n200 131.29e-18 M=1
c1585 a4 n192 131.29e-18 M=1
c1586 a3 n393 46.88e-18 M=1
c1587 a3 n242 46.88e-18 M=1
c1588 a3 n229 46.88e-18 M=1
c1589 a3 n224 46.88e-18 M=1
c1590 a3 n213 83.84e-18 M=1
c1591 a2 n405 46.88e-18 M=1
c1592 a2 n276 131.29e-18 M=1
c1593 a2 n267 131.29e-18 M=1
c1594 a1 n407 46.88e-18 M=1
c1595 a1 n323 46.88e-18 M=1
c1596 a1 n312 46.88e-18 M=1
c1597 a1 n305 46.88e-18 M=1
c1598 a1 n291 83.84e-18 M=1
c1599 a0 n419 46.88e-18 M=1
c1600 a0 n356 131.29e-18 M=1
c1601 a0 n348 131.29e-18 M=1
c1602 b15 n417 46.88e-18 M=1
c1603 b15 n350 131.29e-18 M=1
c1604 b15 n345 131.29e-18 M=1
c1605 b14 n406 46.88e-18 M=1
c1606 b14 n316 46.88e-18 M=1
c1607 b14 n306 46.88e-18 M=1
c1608 b14 n299 46.88e-18 M=1
c1609 b14 n284 83.84e-18 M=1
c1610 b13 n403 46.88e-18 M=1
c1611 b13 n268 131.29e-18 M=1
c1612 b13 n261 131.29e-18 M=1
c1613 b12 n392 46.88e-18 M=1
c1614 b12 n235 46.88e-18 M=1
c1615 b12 n226 46.88e-18 M=1
c1616 b12 n218 46.88e-18 M=1
c1617 b12 n209 83.84e-18 M=1
c1618 b11 n389 46.88e-18 M=1
c1619 b11 n194 131.29e-18 M=1
c1620 b11 n189 131.29e-18 M=1
c1621 b10 n378 46.88e-18 M=1
c1622 b10 n160 46.88e-18 M=1
c1623 b10 n150 46.88e-18 M=1
c1624 b10 n143 46.88e-18 M=1
c1625 b10 n128 83.84e-18 M=1
c1626 gnd n358 1.11344e-15 M=1
c1627 gnd n357 341.44e-18 M=1
c1628 gnd n356 354.4e-18 M=1
c1629 gnd n354 874.5e-18 M=1
c1630 gnd n350 354.4e-18 M=1
c1631 gnd n349 771.36e-18 M=1
c1632 gnd n348 585.12e-18 M=1
c1633 gnd n346 83.72e-18 M=1
c1634 gnd n345 585.12e-18 M=1
c1635 gnd n344 354.4e-18 M=1
c1636 gnd n343 611.2e-18 M=1
c1637 gnd n342 220.32e-18 M=1
c1638 gnd n340 585.12e-18 M=1
c1639 gnd n338 129.58e-18 M=1
c1640 gnd n337 195e-18 M=1
c1641 gnd n335 195e-18 M=1
c1642 gnd n333 354.4e-18 M=1
c1643 gnd n331 129.58e-18 M=1
c1644 gnd n328 171.98e-18 M=1
c1645 gnd n327 611.2e-18 M=1
c1646 gnd n323 129.58e-18 M=1
c1647 gnd n321 354.4e-18 M=1
c1648 gnd n318 771.36e-18 M=1
c1649 gnd n317 771.36e-18 M=1
c1650 gnd n316 129.58e-18 M=1
c1651 gnd n315 585.12e-18 M=1
c1652 gnd n313 585.12e-18 M=1
c1653 gnd n312 585.12e-18 M=1
c1654 gnd n311 611.2e-18 M=1
c1655 gnd n310 124.5e-18 M=1
c1656 gnd n307 354.4e-18 M=1
c1657 gnd n306 585.12e-18 M=1
c1658 gnd n305 354.4e-18 M=1
c1659 gnd n304 195e-18 M=1
c1660 gnd n303 195e-18 M=1
c1661 gnd n299 354.4e-18 M=1
c1662 gnd n298 124.5e-18 M=1
c1663 gnd n297 611.2e-18 M=1
c1664 gnd n296 354.4e-18 M=1
c1665 gnd n291 985.56e-18 M=1
c1666 gnd n290 771.36e-18 M=1
c1667 gnd n289 585.12e-18 M=1
c1668 gnd n286 585.12e-18 M=1
c1669 gnd n285 771.36e-18 M=1
c1670 gnd n284 757.6e-18 M=1
c1671 gnd n281 757.6e-18 M=1
c1672 gnd n279 354.4e-18 M=1
c1673 gnd n278 611.2e-18 M=1
c1674 gnd n277 124.5e-18 M=1
c1675 gnd n276 354.4e-18 M=1
c1676 gnd n272 985.56e-18 M=1
c1677 gnd n270 195e-18 M=1
c1678 gnd n269 195e-18 M=1
c1679 gnd n268 354.4e-18 M=1
c1680 gnd n267 585.12e-18 M=1
c1681 gnd n266 354.4e-18 M=1
c1682 gnd n264 124.5e-18 M=1
c1683 gnd n263 611.2e-18 M=1
c1684 gnd n261 585.12e-18 M=1
c1685 gnd n260 585.12e-18 M=1
c1686 gnd n258 585.12e-18 M=1
c1687 gnd n257 129.58e-18 M=1
c1688 gnd n256 771.36e-18 M=1
c1689 gnd n255 771.36e-18 M=1
c1690 gnd n252 354.4e-18 M=1
c1691 gnd n250 129.58e-18 M=1
c1692 gnd n247 611.2e-18 M=1
c1693 gnd n246 171.98e-18 M=1
c1694 gnd n242 129.58e-18 M=1
c1695 gnd n240 354.4e-18 M=1
c1696 gnd n238 195e-18 M=1
c1697 gnd n236 195e-18 M=1
c1698 gnd n235 129.58e-18 M=1
c1699 gnd n234 585.12e-18 M=1
c1700 gnd n232 220.32e-18 M=1
c1701 gnd n231 611.2e-18 M=1
c1702 gnd n230 354.4e-18 M=1
c1703 gnd n229 585.12e-18 M=1
c1704 gnd n226 585.12e-18 M=1
c1705 gnd n225 771.36e-18 M=1
c1706 gnd n224 354.4e-18 M=1
c1707 gnd n220 83.72e-18 M=1
c1708 gnd n218 354.4e-18 M=1
c1709 gnd n217 341.44e-18 M=1
c1710 gnd n215 1.56886e-15 M=1
c1711 gnd n213 874.5e-18 M=1
c1712 gnd n209 1.11344e-15 M=1
c1713 gnd n204 1.56886e-15 M=1
c1714 gnd n202 1.11344e-15 M=1
c1715 gnd n201 341.44e-18 M=1
c1716 gnd n200 354.4e-18 M=1
c1717 gnd n198 874.5e-18 M=1
c1718 gnd n194 354.4e-18 M=1
c1719 gnd n193 771.36e-18 M=1
c1720 gnd n192 585.12e-18 M=1
c1721 gnd n190 83.72e-18 M=1
c1722 gnd n189 585.12e-18 M=1
c1723 gnd n188 354.4e-18 M=1
c1724 gnd n187 611.2e-18 M=1
c1725 gnd n186 220.32e-18 M=1
c1726 gnd n184 585.12e-18 M=1
c1727 gnd n182 129.58e-18 M=1
c1728 gnd n181 195e-18 M=1
c1729 gnd n179 195e-18 M=1
c1730 gnd n177 354.4e-18 M=1
c1731 gnd n175 129.58e-18 M=1
c1732 gnd n172 171.98e-18 M=1
c1733 gnd n171 611.2e-18 M=1
c1734 gnd n167 129.58e-18 M=1
c1735 gnd n165 354.4e-18 M=1
c1736 gnd n162 771.36e-18 M=1
c1737 gnd n161 771.36e-18 M=1
c1738 gnd n160 129.58e-18 M=1
c1739 gnd n159 585.12e-18 M=1
c1740 gnd n157 585.12e-18 M=1
c1741 gnd n156 585.12e-18 M=1
c1742 gnd n155 611.2e-18 M=1
c1743 gnd n154 124.5e-18 M=1
c1744 gnd n151 354.4e-18 M=1
c1745 gnd n150 585.12e-18 M=1
c1746 gnd n149 354.4e-18 M=1
c1747 gnd n148 195e-18 M=1
c1748 gnd n147 195e-18 M=1
c1749 gnd n143 354.4e-18 M=1
c1750 gnd n142 124.5e-18 M=1
c1751 gnd n141 611.2e-18 M=1
c1752 gnd n140 354.4e-18 M=1
c1753 gnd n135 985.56e-18 M=1
c1754 gnd n134 771.36e-18 M=1
c1755 gnd n133 585.12e-18 M=1
c1756 gnd n130 585.12e-18 M=1
c1757 gnd n129 771.36e-18 M=1
c1758 gnd n128 757.6e-18 M=1
c1759 gnd n125 757.6e-18 M=1
c1760 gnd n123 354.4e-18 M=1
c1761 gnd n122 611.2e-18 M=1
c1762 gnd n121 124.5e-18 M=1
c1763 gnd n120 354.4e-18 M=1
c1764 gnd n116 985.56e-18 M=1
c1765 gnd n114 195e-18 M=1
c1766 gnd n113 195e-18 M=1
c1767 gnd n112 354.4e-18 M=1
c1768 gnd n111 585.12e-18 M=1
c1769 gnd n110 354.4e-18 M=1
c1770 gnd n108 124.5e-18 M=1
c1771 gnd n107 611.2e-18 M=1
c1772 gnd n105 585.12e-18 M=1
c1773 gnd n104 585.12e-18 M=1
c1774 gnd n102 585.12e-18 M=1
c1775 gnd n101 129.58e-18 M=1
c1776 gnd n100 771.36e-18 M=1
c1777 gnd n99 771.36e-18 M=1
c1778 gnd n96 354.4e-18 M=1
c1779 gnd n94 129.58e-18 M=1
c1780 gnd n91 611.2e-18 M=1
c1781 gnd n90 171.98e-18 M=1
c1782 gnd n86 129.58e-18 M=1
c1783 gnd n84 354.4e-18 M=1
c1784 gnd n82 195e-18 M=1
c1785 gnd n80 195e-18 M=1
c1786 gnd n79 129.58e-18 M=1
c1787 gnd n78 585.12e-18 M=1
c1788 gnd n76 220.32e-18 M=1
c1789 gnd n75 611.2e-18 M=1
c1790 gnd n74 354.4e-18 M=1
c1791 gnd n73 585.12e-18 M=1
c1792 gnd n70 585.12e-18 M=1
c1793 gnd n69 771.36e-18 M=1
c1794 gnd n68 354.4e-18 M=1
c1795 gnd n64 83.72e-18 M=1
c1796 gnd n62 354.4e-18 M=1
c1797 gnd n61 341.44e-18 M=1
c1798 gnd n59 480.7e-18 M=1
c1799 gnd n57 874.5e-18 M=1
c1800 gnd n53 1.11344e-15 M=1
c1801 gnd a9 942.4e-18 M=1
c1802 gnd a8 129.4e-18 M=1
c1803 gnd a7 942.4e-18 M=1
c1804 gnd a6 129.4e-18 M=1
c1805 gnd a5 942.4e-18 M=1
c1806 gnd a4 129.4e-18 M=1
c1807 gnd a3 942.4e-18 M=1
c1808 gnd a2 129.4e-18 M=1
c1809 gnd a1 942.4e-18 M=1
c1810 gnd a0 129.4e-18 M=1
c1811 gnd b15 129.4e-18 M=1
c1812 gnd b14 942.4e-18 M=1
c1813 gnd b13 129.4e-18 M=1
c1814 gnd b12 942.4e-18 M=1
c1815 gnd b11 129.4e-18 M=1
c1816 gnd b10 942.4e-18 M=1
c1817 a15 n417 46.88e-18 M=1
c1818 a15 n354 83.84e-18 M=1
c1819 a15 n350 46.88e-18 M=1
c1820 a15 n345 46.88e-18 M=1
c1821 a15 n331 46.88e-18 M=1
c1822 a15 b15 140.64e-18 M=1
c1823 a15 gnd 942.4e-18 M=1
c1824 a14 n406 46.88e-18 M=1
c1825 a14 n306 131.29e-18 M=1
c1826 a14 n299 131.29e-18 M=1
c1827 a14 b14 140.64e-18 M=1
c1828 a14 gnd 129.4e-18 M=1
c1829 a13 n403 46.88e-18 M=1
c1830 a13 n272 83.84e-18 M=1
c1831 a13 n268 46.88e-18 M=1
c1832 a13 n261 46.88e-18 M=1
c1833 a13 n250 46.88e-18 M=1
c1834 a13 b13 140.64e-18 M=1
c1835 a13 gnd 942.4e-18 M=1
c1836 a12 n392 46.88e-18 M=1
c1837 a12 n226 131.29e-18 M=1
c1838 a12 n218 131.29e-18 M=1
c1839 a12 b12 140.64e-18 M=1
c1840 a12 gnd 129.4e-18 M=1
c1841 a11 n389 46.88e-18 M=1
c1842 a11 n198 83.84e-18 M=1
c1843 a11 n194 46.88e-18 M=1
c1844 a11 n189 46.88e-18 M=1
c1845 a11 n175 46.88e-18 M=1
c1846 a11 b11 140.64e-18 M=1
c1847 a11 gnd 942.4e-18 M=1
c1848 a10 n378 46.88e-18 M=1
c1849 a10 n150 131.29e-18 M=1
c1850 a10 n143 131.29e-18 M=1
c1851 a10 b10 140.64e-18 M=1
c1852 a10 gnd 129.4e-18 M=1
c1853 cin n412 46.88e-18 M=1
c1854 cin n395 46.88e-18 M=1
c1855 cin n358 93.76e-18 M=1
c1856 cin n349 84.6e-18 M=1
c1857 cin n343 84.6e-18 M=1
c1858 cin n340 46.88e-18 M=1
c1859 cin n333 131.29e-18 M=1
c1860 cin n332 46.88e-18 M=1
c1861 cin n232 46.88e-18 M=1
c1862 cin n230 46.88e-18 M=1
c1863 cin n217 46.88e-18 M=1
c1864 cin gnd 659.295e-18 M=1
c1865 s15 n413 85.36e-18 M=1
c1866 s15 n354 83.84e-18 M=1
c1867 s15 n321 83.84e-18 M=1
c1868 s15 n315 83.84e-18 M=1
c1869 s14 n410 85.36e-18 M=1
c1870 s14 n296 83.84e-18 M=1
c1871 s14 n289 83.84e-18 M=1
c1872 s14 n284 83.84e-18 M=1
c1873 s13 n402 85.36e-18 M=1
c1874 s13 n272 83.84e-18 M=1
c1875 s13 n266 83.84e-18 M=1
c1876 s13 n260 83.84e-18 M=1
c1877 s12 n398 85.36e-18 M=1
c1878 s12 n240 83.84e-18 M=1
c1879 s12 n234 83.84e-18 M=1
c1880 s12 n209 83.84e-18 M=1
c1881 s11 n385 85.36e-18 M=1
c1882 s11 n198 83.84e-18 M=1
c1883 s11 n165 83.84e-18 M=1
c1884 s11 n159 83.84e-18 M=1
c1885 s10 n382 85.36e-18 M=1
c1886 s10 n140 83.84e-18 M=1
c1887 s10 n133 83.84e-18 M=1
c1888 s10 n128 83.84e-18 M=1
c1889 cout gnd 599.36e-18 M=1
c1890 b9 n375 46.88e-18 M=1
c1891 b9 n112 131.29e-18 M=1
c1892 b9 n105 131.29e-18 M=1
c1893 b9 a9 140.64e-18 M=1
c1894 b9 gnd 129.4e-18 M=1
c1895 b8 n364 46.88e-18 M=1
c1896 b8 n79 46.88e-18 M=1
c1897 b8 n70 46.88e-18 M=1
c1898 b8 n62 46.88e-18 M=1
c1899 b8 n53 83.84e-18 M=1
c1900 b8 a8 140.64e-18 M=1
c1901 b8 gnd 942.4e-18 M=1
c1902 b7 n365 46.88e-18 M=1
c1903 b7 n73 131.29e-18 M=1
c1904 b7 n68 131.29e-18 M=1
c1905 b7 a7 140.64e-18 M=1
c1906 b7 gnd 129.4e-18 M=1
c1907 b6 n377 46.88e-18 M=1
c1908 b6 n125 83.84e-18 M=1
c1909 b6 n120 46.88e-18 M=1
c1910 b6 n111 46.88e-18 M=1
c1911 b6 n101 46.88e-18 M=1
c1912 b6 a6 140.64e-18 M=1
c1913 b6 gnd 942.4e-18 M=1
c1914 b5 n379 46.88e-18 M=1
c1915 b5 n156 131.29e-18 M=1
c1916 b5 n149 131.29e-18 M=1
c1917 b5 a5 140.64e-18 M=1
c1918 b5 gnd 129.4e-18 M=1
c1919 b4 n391 46.88e-18 M=1
c1920 b4 n202 83.84e-18 M=1
c1921 b4 n200 46.88e-18 M=1
c1922 b4 n192 46.88e-18 M=1
c1923 b4 n182 46.88e-18 M=1
c1924 b4 a4 140.64e-18 M=1
c1925 b4 gnd 942.4e-18 M=1
c1926 s9 n374 85.36e-18 M=1
c1927 s9 n116 83.84e-18 M=1
c1928 s9 n110 83.84e-18 M=1
c1929 s9 n104 83.84e-18 M=1
c1930 b3 n393 46.88e-18 M=1
c1931 b3 n229 131.29e-18 M=1
c1932 b3 n224 131.29e-18 M=1
c1933 b3 a3 140.64e-18 M=1
c1934 b3 gnd 129.4e-18 M=1
c1935 s8 n370 85.36e-18 M=1
c1936 s8 n84 83.84e-18 M=1
c1937 s8 n78 83.84e-18 M=1
c1938 s8 n53 83.84e-18 M=1
c1939 b2 n405 46.88e-18 M=1
c1940 b2 n281 83.84e-18 M=1
c1941 b2 n276 46.88e-18 M=1
c1942 b2 n267 46.88e-18 M=1
c1943 b2 n257 46.88e-18 M=1
c1944 b2 a2 140.64e-18 M=1
c1945 b2 gnd 942.4e-18 M=1
c1946 s7 n369 85.36e-18 M=1
c1947 s7 n102 83.84e-18 M=1
c1948 s7 n96 83.84e-18 M=1
c1949 s7 n57 83.84e-18 M=1
c1950 b1 n407 46.88e-18 M=1
c1951 b1 n312 131.29e-18 M=1
c1952 b1 n305 131.29e-18 M=1
c1953 b1 a1 140.64e-18 M=1
c1954 b1 gnd 129.4e-18 M=1
c1955 s6 n373 85.36e-18 M=1
c1956 s6 n130 83.84e-18 M=1
c1957 s6 n125 83.84e-18 M=1
c1958 s6 n123 83.84e-18 M=1
c1959 b0 n419 46.88e-18 M=1
c1960 b0 n358 83.84e-18 M=1
c1961 b0 n356 46.88e-18 M=1
c1962 b0 n348 46.88e-18 M=1
c1963 b0 n338 46.88e-18 M=1
c1964 b0 a0 140.64e-18 M=1
c1965 b0 gnd 942.4e-18 M=1
c1966 s5 n380 85.36e-18 M=1
c1967 s5 n157 83.84e-18 M=1
c1968 s5 n151 83.84e-18 M=1
c1969 s5 n135 83.84e-18 M=1
c1970 vdd n435 346.18e-18 M=1
c1971 vdd n434 631.26e-18 M=1
c1972 vdd n433 631.26e-18 M=1
c1973 vdd n432 631.26e-18 M=1
c1974 vdd n431 631.26e-18 M=1
c1975 vdd n430 631.26e-18 M=1
c1976 vdd n429 631.26e-18 M=1
c1977 vdd n428 346.18e-18 M=1
c1978 vdd n427 346.18e-18 M=1
c1979 vdd n426 631.26e-18 M=1
c1980 vdd n425 631.26e-18 M=1
c1981 vdd n424 631.26e-18 M=1
c1982 vdd n423 631.26e-18 M=1
c1983 vdd n422 631.26e-18 M=1
c1984 vdd n421 631.26e-18 M=1
c1985 vdd n420 346.18e-18 M=1
c1986 vdd n419 85.36e-18 M=1
c1987 vdd n417 85.36e-18 M=1
c1988 vdd n416 85.36e-18 M=1
c1989 vdd n413 85.36e-18 M=1
c1990 vdd n412 85.36e-18 M=1
c1991 vdd n410 85.36e-18 M=1
c1992 vdd n408 85.36e-18 M=1
c1993 vdd n407 85.36e-18 M=1
c1994 vdd n406 85.36e-18 M=1
c1995 vdd n405 85.36e-18 M=1
c1996 vdd n403 85.36e-18 M=1
c1997 vdd n402 85.36e-18 M=1
c1998 vdd n401 85.36e-18 M=1
c1999 vdd n398 85.36e-18 M=1
c2000 vdd n397 85.36e-18 M=1
c2001 vdd n395 85.36e-18 M=1
c2002 vdd n393 85.36e-18 M=1
c2003 vdd n392 85.36e-18 M=1
c2004 vdd n391 85.36e-18 M=1
c2005 vdd n389 85.36e-18 M=1
c2006 vdd n388 85.36e-18 M=1
c2007 vdd n385 85.36e-18 M=1
c2008 vdd n384 85.36e-18 M=1
c2009 vdd n382 85.36e-18 M=1
c2010 vdd n380 85.36e-18 M=1
c2011 vdd n379 85.36e-18 M=1
c2012 vdd n378 85.36e-18 M=1
c2013 vdd n377 85.36e-18 M=1
c2014 vdd n375 85.36e-18 M=1
c2015 vdd n374 85.36e-18 M=1
c2016 vdd n373 85.36e-18 M=1
c2017 vdd n370 85.36e-18 M=1
c2018 vdd n369 85.36e-18 M=1
c2019 vdd n367 85.36e-18 M=1
c2020 vdd n365 85.36e-18 M=1
c2021 vdd n364 85.36e-18 M=1
c2022 vdd n358 47.84e-18 M=1
c2023 vdd n357 548.93e-18 M=1
c2024 vdd n356 83.36e-18 M=1
c2025 vdd n354 167.98e-18 M=1
c2026 vdd n350 83.36e-18 M=1
c2027 vdd n348 47.84e-18 M=1
c2028 vdd n346 95.32e-18 M=1
c2029 vdd n345 47.84e-18 M=1
c2030 vdd n344 83.36e-18 M=1
c2031 vdd n340 47.84e-18 M=1
c2032 vdd n338 133.54e-18 M=1
c2033 vdd n337 199.32e-18 M=1
c2034 vdd n335 199.32e-18 M=1
c2035 vdd n333 83.36e-18 M=1
c2036 vdd n331 133.54e-18 M=1
c2037 vdd n328 969.21e-18 M=1
c2038 vdd n323 133.54e-18 M=1
c2039 vdd n321 83.36e-18 M=1
c2040 vdd n316 133.54e-18 M=1
c2041 vdd n315 47.84e-18 M=1
c2042 vdd n313 47.84e-18 M=1
c2043 vdd n312 47.84e-18 M=1
c2044 vdd n310 836.93e-18 M=1
c2045 vdd n307 83.36e-18 M=1
c2046 vdd n306 47.84e-18 M=1
c2047 vdd n305 83.36e-18 M=1
c2048 vdd n304 199.32e-18 M=1
c2049 vdd n303 199.32e-18 M=1
c2050 vdd n299 83.36e-18 M=1
c2051 vdd n298 836.93e-18 M=1
c2052 vdd n296 83.36e-18 M=1
c2053 vdd n291 130.84e-18 M=1
c2054 vdd n289 47.84e-18 M=1
c2055 vdd n286 47.84e-18 M=1
c2056 vdd n279 83.36e-18 M=1
c2057 vdd n277 836.93e-18 M=1
c2058 vdd n276 83.36e-18 M=1
c2059 vdd n272 130.84e-18 M=1
c2060 vdd n270 199.32e-18 M=1
c2061 vdd n269 199.32e-18 M=1
c2062 vdd n268 83.36e-18 M=1
c2063 vdd n267 47.84e-18 M=1
c2064 vdd n266 83.36e-18 M=1
c2065 vdd n264 836.93e-18 M=1
c2066 vdd n261 47.84e-18 M=1
c2067 vdd n260 47.84e-18 M=1
c2068 vdd n258 47.84e-18 M=1
c2069 vdd n257 133.54e-18 M=1
c2070 vdd n252 83.36e-18 M=1
c2071 vdd n250 133.54e-18 M=1
c2072 vdd n246 969.21e-18 M=1
c2073 vdd n242 133.54e-18 M=1
c2074 vdd n240 83.36e-18 M=1
c2075 vdd n238 199.32e-18 M=1
c2076 vdd n236 199.32e-18 M=1
c2077 vdd n235 133.54e-18 M=1
c2078 vdd n234 47.84e-18 M=1
c2079 vdd n230 83.36e-18 M=1
c2080 vdd n229 47.84e-18 M=1
c2081 vdd n226 47.84e-18 M=1
c2082 vdd n224 83.36e-18 M=1
c2083 vdd n220 95.32e-18 M=1
c2084 vdd n218 83.36e-18 M=1
c2085 vdd n217 548.93e-18 M=1
c2086 vdd n215 1.11167e-15 M=1
c2087 vdd n213 167.98e-18 M=1
c2088 vdd n209 47.84e-18 M=1
c2089 vdd n204 1.11167e-15 M=1
c2090 vdd n202 47.84e-18 M=1
c2091 vdd n201 548.93e-18 M=1
c2092 vdd n200 83.36e-18 M=1
c2093 vdd n198 167.98e-18 M=1
c2094 vdd n194 83.36e-18 M=1
c2095 vdd n192 47.84e-18 M=1
c2096 vdd n190 95.32e-18 M=1
c2097 vdd n189 47.84e-18 M=1
c2098 vdd n188 83.36e-18 M=1
c2099 vdd n184 47.84e-18 M=1
c2100 vdd n182 133.54e-18 M=1
c2101 vdd n181 199.32e-18 M=1
c2102 vdd n179 199.32e-18 M=1
c2103 vdd n177 83.36e-18 M=1
c2104 vdd n175 133.54e-18 M=1
c2105 vdd n172 969.21e-18 M=1
c2106 vdd n167 133.54e-18 M=1
c2107 vdd n165 83.36e-18 M=1
c2108 vdd n160 133.54e-18 M=1
c2109 vdd n159 47.84e-18 M=1
c2110 vdd n157 47.84e-18 M=1
c2111 vdd n156 47.84e-18 M=1
c2112 vdd n154 836.93e-18 M=1
c2113 vdd n151 83.36e-18 M=1
c2114 vdd n150 47.84e-18 M=1
c2115 vdd n149 83.36e-18 M=1
c2116 vdd n148 199.32e-18 M=1
c2117 vdd n147 199.32e-18 M=1
c2118 vdd n143 83.36e-18 M=1
c2119 vdd n142 836.93e-18 M=1
c2120 vdd n140 83.36e-18 M=1
c2121 vdd n135 130.84e-18 M=1
c2122 vdd n133 47.84e-18 M=1
c2123 vdd n130 47.84e-18 M=1
c2124 vdd n123 83.36e-18 M=1
c2125 vdd n121 836.93e-18 M=1
c2126 vdd n120 83.36e-18 M=1
c2127 vdd n116 130.84e-18 M=1
c2128 vdd n114 199.32e-18 M=1
c2129 vdd n113 199.32e-18 M=1
c2130 vdd n112 83.36e-18 M=1
c2131 vdd n111 47.84e-18 M=1
c2132 vdd n110 83.36e-18 M=1
c2133 vdd n108 836.93e-18 M=1
c2134 vdd n105 47.84e-18 M=1
c2135 vdd n104 47.84e-18 M=1
c2136 vdd n102 47.84e-18 M=1
c2137 vdd n101 133.54e-18 M=1
c2138 vdd n96 83.36e-18 M=1
c2139 vdd n94 133.54e-18 M=1
c2140 vdd n90 969.21e-18 M=1
c2141 vdd n86 133.54e-18 M=1
c2142 vdd n84 83.36e-18 M=1
c2143 vdd n82 199.32e-18 M=1
c2144 vdd n80 199.32e-18 M=1
c2145 vdd n79 133.54e-18 M=1
c2146 vdd n78 47.84e-18 M=1
c2147 vdd n74 83.36e-18 M=1
c2148 vdd n73 47.84e-18 M=1
c2149 vdd n70 47.84e-18 M=1
c2150 vdd n68 83.36e-18 M=1
c2151 vdd n64 95.32e-18 M=1
c2152 vdd n62 83.36e-18 M=1
c2153 vdd n61 548.93e-18 M=1
c2154 vdd n59 1.02831e-15 M=1
c2155 vdd n57 167.98e-18 M=1
c2156 vdd n53 47.84e-18 M=1
c2157 vdd a9 67e-18 M=1
c2158 vdd a8 679.86e-18 M=1
c2159 vdd a7 67e-18 M=1
c2160 vdd a6 679.86e-18 M=1
c2161 vdd a5 67e-18 M=1
c2162 vdd a4 679.86e-18 M=1
c2163 vdd a3 67e-18 M=1
c2164 vdd a2 679.86e-18 M=1
c2165 vdd a1 67e-18 M=1
c2166 vdd a0 679.86e-18 M=1
c2167 vdd b15 679.86e-18 M=1
c2168 vdd b14 67e-18 M=1
c2169 vdd b13 679.86e-18 M=1
c2170 vdd b12 67e-18 M=1
c2171 vdd b11 679.86e-18 M=1
c2172 vdd b10 67e-18 M=1
c2173 vdd gnd 47.4713e-15 M=1
c2174 vdd a15 67e-18 M=1
c2175 vdd a14 679.86e-18 M=1
c2176 vdd a13 67e-18 M=1
c2177 vdd a12 679.86e-18 M=1
c2178 vdd a11 67e-18 M=1
c2179 vdd a10 679.86e-18 M=1
c2180 vdd cin 1.02831e-15 M=1
c2181 vdd cout 301.12e-18 M=1
c2182 vdd b9 679.86e-18 M=1
c2183 vdd b8 67e-18 M=1
c2184 vdd b7 679.86e-18 M=1
c2185 vdd b6 67e-18 M=1
c2186 vdd b5 679.86e-18 M=1
c2187 vdd b4 67e-18 M=1
c2188 vdd b3 679.86e-18 M=1
c2189 vdd b2 67e-18 M=1
c2190 vdd b1 679.86e-18 M=1
c2191 vdd b0 67e-18 M=1
c2192 s4 n384 85.36e-18 M=1
c2193 s4 n202 83.84e-18 M=1
c2194 s4 n184 83.84e-18 M=1
c2195 s4 n177 83.84e-18 M=1
c2196 s3 n397 85.36e-18 M=1
c2197 s3 n258 83.84e-18 M=1
c2198 s3 n252 83.84e-18 M=1
c2199 s3 n213 83.84e-18 M=1
c2200 n354 n363 49.16e-18 M=1
c2201 n342 n357 79.36e-18 M=1
c2202 n342 n344 79.36e-18 M=1
c2203 n332 n349 79.36e-18 M=1
c2204 n318 n324 79.36e-18 M=1
c2205 n317 n330 79.36e-18 M=1
c2206 n310 n354 194.48e-18 M=1
c2207 n310 n318 35.365e-18 M=1
c2208 n297 n354 47.44e-18 M=1
c2209 n291 n328 79.36e-18 M=1
c2210 n291 n317 165.055e-18 M=1
c2211 n290 n322 79.36e-18 M=1
c2212 n281 n298 79.36e-18 M=1
c2213 n277 n284 79.36e-18 M=1
c2214 n272 n351 49.16e-18 M=1
c2215 n256 n272 165.055e-18 M=1
c2216 n255 n264 35.365e-18 M=1
c2217 n251 n285 79.36e-18 M=1
c2218 n249 n255 79.36e-18 M=1
c2219 n246 n272 79.36e-18 M=1
c2220 n244 n256 79.36e-18 M=1
c2221 n230 n232 79.36e-18 M=1
c2222 n225 n241 79.36e-18 M=1
c2223 n223 n291 49.16e-18 M=1
c2224 n217 n232 79.36e-18 M=1
c2225 n213 n278 47.44e-18 M=1
c2226 n213 n264 194.48e-18 M=1
c2227 n210 n213 49.16e-18 M=1
c2228 n204 n234 219.98e-18 M=1
c2229 n204 n209 158.72e-18 M=1
c2230 n202 n215 158.72e-18 M=1
c2231 n198 n208 49.16e-18 M=1
c2232 n186 n201 79.36e-18 M=1
c2233 n186 n188 79.36e-18 M=1
c2234 n184 n215 219.98e-18 M=1
c2235 n176 n193 79.36e-18 M=1
c2236 n162 n168 79.36e-18 M=1
c2237 n161 n174 79.36e-18 M=1
c2238 n154 n198 194.48e-18 M=1
c2239 n154 n162 35.365e-18 M=1
c2240 n141 n198 47.44e-18 M=1
c2241 n135 n172 79.36e-18 M=1
c2242 n135 n161 165.055e-18 M=1
c2243 n134 n166 79.36e-18 M=1
c2244 n125 n142 79.36e-18 M=1
c2245 n121 n128 79.36e-18 M=1
c2246 n116 n195 49.16e-18 M=1
c2247 n100 n116 165.055e-18 M=1
c2248 n99 n108 35.365e-18 M=1
c2249 n95 n129 79.36e-18 M=1
c2250 n93 n99 79.36e-18 M=1
c2251 n90 n116 79.36e-18 M=1
c2252 n88 n100 79.36e-18 M=1
c2253 n74 n76 79.36e-18 M=1
c2254 n69 n85 79.36e-18 M=1
c2255 n67 n135 49.16e-18 M=1
c2256 n61 n76 79.36e-18 M=1
c2257 n59 n78 219.98e-18 M=1
c2258 n57 n122 47.44e-18 M=1
c2259 n57 n108 194.48e-18 M=1
c2260 n54 n57 49.16e-18 M=1
c2261 n53 n59 158.72e-18 M=1
c2262 gnd n358 1.543e-15 M=1
c2263 gnd n354 985.11e-18 M=1
c2264 gnd n342 144.56e-18 M=1
c2265 gnd n332 870.26e-18 M=1
c2266 gnd n330 866.18e-18 M=1
c2267 gnd n324 754.49e-18 M=1
c2268 gnd n322 856.1e-18 M=1
c2269 gnd n291 1.28234e-15 M=1
c2270 gnd n284 1.35108e-15 M=1
c2271 gnd n281 1.35108e-15 M=1
c2272 gnd n272 1.28234e-15 M=1
c2273 gnd n251 856.1e-18 M=1
c2274 gnd n249 754.49e-18 M=1
c2275 gnd n244 866.18e-18 M=1
c2276 gnd n241 870.26e-18 M=1
c2277 gnd n232 144.56e-18 M=1
c2278 gnd n215 420.74e-18 M=1
c2279 gnd n213 985.11e-18 M=1
c2280 gnd n209 1.543e-15 M=1
c2281 gnd n204 420.74e-18 M=1
c2282 gnd n202 1.543e-15 M=1
c2283 gnd n198 985.11e-18 M=1
c2284 gnd n186 144.56e-18 M=1
c2285 gnd n176 870.26e-18 M=1
c2286 gnd n174 866.18e-18 M=1
c2287 gnd n168 754.49e-18 M=1
c2288 gnd n166 856.1e-18 M=1
c2289 gnd n135 1.28234e-15 M=1
c2290 gnd n128 1.35108e-15 M=1
c2291 gnd n125 1.35108e-15 M=1
c2292 gnd n116 1.28234e-15 M=1
c2293 gnd n95 856.1e-18 M=1
c2294 gnd n93 754.49e-18 M=1
c2295 gnd n88 866.18e-18 M=1
c2296 gnd n85 870.26e-18 M=1
c2297 gnd n76 144.56e-18 M=1
c2298 gnd n59 1.2269e-15 M=1
c2299 gnd n57 985.11e-18 M=1
c2300 gnd n53 1.543e-15 M=1
c2301 gnd a9 92.31e-18 M=1
c2302 gnd a8 60.12e-18 M=1
c2303 gnd a7 92.31e-18 M=1
c2304 gnd a6 60.12e-18 M=1
c2305 gnd a5 92.31e-18 M=1
c2306 gnd a4 60.12e-18 M=1
c2307 gnd a3 92.31e-18 M=1
c2308 gnd a2 60.12e-18 M=1
c2309 gnd a1 92.31e-18 M=1
c2310 gnd a0 60.12e-18 M=1
c2311 gnd b15 60.12e-18 M=1
c2312 gnd b14 92.31e-18 M=1
c2313 gnd b13 65.68e-18 M=1
c2314 gnd b12 100.747e-18 M=1
c2315 gnd b11 60.12e-18 M=1
c2316 gnd b10 92.31e-18 M=1
c2317 a15 b15 79.36e-18 M=1
c2318 a15 gnd 92.31e-18 M=1
c2319 a14 b14 79.36e-18 M=1
c2320 a14 gnd 65.6475e-18 M=1
c2321 a13 b13 79.36e-18 M=1
c2322 a13 gnd 92.31e-18 M=1
c2323 a12 b12 79.36e-18 M=1
c2324 a12 gnd 60.12e-18 M=1
c2325 a11 b11 79.36e-18 M=1
c2326 a11 gnd 92.31e-18 M=1
c2327 a10 b10 79.36e-18 M=1
c2328 a10 gnd 60.12e-18 M=1
c2329 cin n358 158.72e-18 M=1
c2330 cin n340 219.98e-18 M=1
c2331 cin gnd 103.82e-18 M=1
c2332 b9 a9 79.36e-18 M=1
c2333 b9 gnd 60.12e-18 M=1
c2334 b8 a8 79.36e-18 M=1
c2335 b8 gnd 97.8375e-18 M=1
c2336 b7 a7 79.36e-18 M=1
c2337 b7 gnd 60.12e-18 M=1
c2338 b6 a6 79.36e-18 M=1
c2339 b6 gnd 92.31e-18 M=1
c2340 b5 a5 79.36e-18 M=1
c2341 b5 gnd 60.12e-18 M=1
c2342 b4 a4 79.36e-18 M=1
c2343 b4 gnd 92.31e-18 M=1
c2344 b3 a3 79.36e-18 M=1
c2345 b3 gnd 62.965e-18 M=1
c2346 b2 a2 79.36e-18 M=1
c2347 b2 gnd 92.31e-18 M=1
c2348 b1 a1 79.36e-18 M=1
c2349 b1 gnd 60.12e-18 M=1
c2350 b0 a0 79.36e-18 M=1
c2351 b0 gnd 92.31e-18 M=1
c2352 vdd n358 320.3e-18 M=1
c2353 vdd n357 418.32e-18 M=1
c2354 vdd n354 519.35e-18 M=1
c2355 vdd n342 418.32e-18 M=1
c2356 vdd n328 532.06e-18 M=1
c2357 vdd n324 21.46e-18 M=1
c2358 vdd n310 478.785e-18 M=1
c2359 vdd n298 491.4e-18 M=1
c2360 vdd n291 536.235e-18 M=1
c2361 vdd n284 606.35e-18 M=1
c2362 vdd n281 606.35e-18 M=1
c2363 vdd n277 491.4e-18 M=1
c2364 vdd n272 536.235e-18 M=1
c2365 vdd n264 478.785e-18 M=1
c2366 vdd n249 21.46e-18 M=1
c2367 vdd n246 532.06e-18 M=1
c2368 vdd n232 418.32e-18 M=1
c2369 vdd n217 418.32e-18 M=1
c2370 vdd n215 743.66e-18 M=1
c2371 vdd n213 519.35e-18 M=1
c2372 vdd n209 320.3e-18 M=1
c2373 vdd n204 743.66e-18 M=1
c2374 vdd n202 320.3e-18 M=1
c2375 vdd n201 418.32e-18 M=1
c2376 vdd n198 519.35e-18 M=1
c2377 vdd n186 418.32e-18 M=1
c2378 vdd n172 532.06e-18 M=1
c2379 vdd n168 21.46e-18 M=1
c2380 vdd n154 478.785e-18 M=1
c2381 vdd n142 491.4e-18 M=1
c2382 vdd n135 536.235e-18 M=1
c2383 vdd n128 606.35e-18 M=1
c2384 vdd n125 606.35e-18 M=1
c2385 vdd n121 491.4e-18 M=1
c2386 vdd n116 536.235e-18 M=1
c2387 vdd n108 478.785e-18 M=1
c2388 vdd n93 21.46e-18 M=1
c2389 vdd n90 532.06e-18 M=1
c2390 vdd n76 418.32e-18 M=1
c2391 vdd n61 418.32e-18 M=1
c2392 vdd n59 743.66e-18 M=1
c2393 vdd n57 519.35e-18 M=1
c2394 vdd n53 320.3e-18 M=1
c2395 vdd a9 390.13e-18 M=1
c2396 vdd a8 357.16e-18 M=1
c2397 vdd a7 390.13e-18 M=1
c2398 vdd a6 357.16e-18 M=1
c2399 vdd a5 390.13e-18 M=1
c2400 vdd a4 357.16e-18 M=1
c2401 vdd a3 390.13e-18 M=1
c2402 vdd a2 357.16e-18 M=1
c2403 vdd a1 390.13e-18 M=1
c2404 vdd a0 357.16e-18 M=1
c2405 vdd b15 357.16e-18 M=1
c2406 vdd b14 390.13e-18 M=1
c2407 vdd b13 357.16e-18 M=1
c2408 vdd b12 394.82e-18 M=1
c2409 vdd b11 357.16e-18 M=1
c2410 vdd b10 390.13e-18 M=1
c2411 vdd a15 390.13e-18 M=1
c2412 vdd a14 357.16e-18 M=1
c2413 vdd a13 390.13e-18 M=1
c2414 vdd a12 357.16e-18 M=1
c2415 vdd a11 390.13e-18 M=1
c2416 vdd a10 357.16e-18 M=1
c2417 vdd cin 536.62e-18 M=1
c2418 vdd b9 357.16e-18 M=1
c2419 vdd b8 390.13e-18 M=1
c2420 vdd b7 357.16e-18 M=1
c2421 vdd b6 390.13e-18 M=1
c2422 vdd b5 357.16e-18 M=1
c2423 vdd b4 390.13e-18 M=1
c2424 vdd b3 362.3e-18 M=1
c2425 vdd b2 390.13e-18 M=1
c2426 vdd b1 357.16e-18 M=1
c2427 vdd b0 390.13e-18 M=1
c2428 n339 n354 191.7e-18 M=1
c2429 n332 n358 88.64e-18 M=1
c2430 n330 n358 88.64e-18 M=1
c2431 n327 n354 23.42e-18 M=1
c2432 n324 n354 88.64e-18 M=1
c2433 n322 n354 177.28e-18 M=1
c2434 n312 n358 28.16e-18 M=1
c2435 n310 n322 56.24e-18 M=1
c2436 n309 n322 83.64e-18 M=1
c2437 n305 n358 28.16e-18 M=1
c2438 n303 n322 28.16e-18 M=1
c2439 n300 n358 56.64e-18 M=1
c2440 n297 n322 28.16e-18 M=1
c2441 n293 n358 56.64e-18 M=1
c2442 n291 n358 233.92e-18 M=1
c2443 n291 n330 88.64e-18 M=1
c2444 n290 n322 28.16e-18 M=1
c2445 n287 n358 56.64e-18 M=1
c2446 n284 n354 88.64e-18 M=1
c2447 n284 n324 88.64e-18 M=1
c2448 n284 n322 88.64e-18 M=1
c2449 n283 n358 56.64e-18 M=1
c2450 n281 n358 233.92e-18 M=1
c2451 n281 n291 177.28e-18 M=1
c2452 n276 n358 28.16e-18 M=1
c2453 n272 n354 88.64e-18 M=1
c2454 n272 n324 88.64e-18 M=1
c2455 n272 n322 88.64e-18 M=1
c2456 n272 n284 177.28e-18 M=1
c2457 n267 n358 28.16e-18 M=1
c2458 n251 n358 88.64e-18 M=1
c2459 n251 n291 88.64e-18 M=1
c2460 n251 n285 28.16e-18 M=1
c2461 n251 n281 88.64e-18 M=1
c2462 n251 n278 28.16e-18 M=1
c2463 n251 n270 28.16e-18 M=1
c2464 n251 n264 56.24e-18 M=1
c2465 n251 n262 83.64e-18 M=1
c2466 n249 n358 88.64e-18 M=1
c2467 n249 n291 88.64e-18 M=1
c2468 n249 n281 88.64e-18 M=1
c2469 n244 n272 88.64e-18 M=1
c2470 n213 n358 88.64e-18 M=1
c2471 n213 n291 88.64e-18 M=1
c2472 n213 n281 88.64e-18 M=1
c2473 n213 n251 177.28e-18 M=1
c2474 n213 n249 88.64e-18 M=1
c2475 n213 n247 23.42e-18 M=1
c2476 n213 n228 191.7e-18 M=1
c2477 n209 n354 88.64e-18 M=1
c2478 n209 n324 88.64e-18 M=1
c2479 n209 n322 88.64e-18 M=1
c2480 n209 n306 28.16e-18 M=1
c2481 n209 n299 28.16e-18 M=1
c2482 n209 n292 56.64e-18 M=1
c2483 n209 n288 56.64e-18 M=1
c2484 n209 n284 233.92e-18 M=1
c2485 n209 n282 56.64e-18 M=1
c2486 n209 n275 56.64e-18 M=1
c2487 n209 n272 233.92e-18 M=1
c2488 n209 n268 28.16e-18 M=1
c2489 n209 n261 28.16e-18 M=1
c2490 n209 n244 88.64e-18 M=1
c2491 n209 n241 88.64e-18 M=1
c2492 n204 n357 28.16e-18 M=1
c2493 n204 n354 649.28e-18 M=1
c2494 n204 n346 55.84e-18 M=1
c2495 n204 n321 28.16e-18 M=1
c2496 n204 n315 28.16e-18 M=1
c2497 n204 n296 28.16e-18 M=1
c2498 n204 n289 28.16e-18 M=1
c2499 n204 n284 677.84e-18 M=1
c2500 n204 n272 725.44e-18 M=1
c2501 n204 n266 28.16e-18 M=1
c2502 n204 n260 28.16e-18 M=1
c2503 n204 n240 28.16e-18 M=1
c2504 n204 n234 28.16e-18 M=1
c2505 n204 n209 408.32e-18 M=1
c2506 n202 n215 408.32e-18 M=1
c2507 n184 n215 28.16e-18 M=1
c2508 n183 n198 191.7e-18 M=1
c2509 n177 n215 28.16e-18 M=1
c2510 n176 n202 88.64e-18 M=1
c2511 n174 n202 88.64e-18 M=1
c2512 n171 n198 23.42e-18 M=1
c2513 n168 n198 88.64e-18 M=1
c2514 n166 n198 177.28e-18 M=1
c2515 n157 n215 28.16e-18 M=1
c2516 n156 n202 28.16e-18 M=1
c2517 n154 n166 56.24e-18 M=1
c2518 n153 n166 83.64e-18 M=1
c2519 n151 n215 28.16e-18 M=1
c2520 n149 n202 28.16e-18 M=1
c2521 n147 n166 28.16e-18 M=1
c2522 n144 n202 56.64e-18 M=1
c2523 n141 n166 28.16e-18 M=1
c2524 n137 n202 56.64e-18 M=1
c2525 n135 n215 725.44e-18 M=1
c2526 n135 n202 233.92e-18 M=1
c2527 n135 n174 88.64e-18 M=1
c2528 n134 n166 28.16e-18 M=1
c2529 n131 n202 56.64e-18 M=1
c2530 n130 n215 28.16e-18 M=1
c2531 n128 n198 88.64e-18 M=1
c2532 n128 n168 88.64e-18 M=1
c2533 n128 n166 88.64e-18 M=1
c2534 n127 n202 56.64e-18 M=1
c2535 n125 n215 677.84e-18 M=1
c2536 n125 n202 233.92e-18 M=1
c2537 n125 n135 177.28e-18 M=1
c2538 n123 n215 28.16e-18 M=1
c2539 n120 n202 28.16e-18 M=1
c2540 n116 n198 88.64e-18 M=1
c2541 n116 n168 88.64e-18 M=1
c2542 n116 n166 88.64e-18 M=1
c2543 n116 n128 177.28e-18 M=1
c2544 n111 n202 28.16e-18 M=1
c2545 n102 n215 28.16e-18 M=1
c2546 n96 n215 28.16e-18 M=1
c2547 n95 n202 88.64e-18 M=1
c2548 n95 n135 88.64e-18 M=1
c2549 n95 n129 28.16e-18 M=1
c2550 n95 n125 88.64e-18 M=1
c2551 n95 n122 28.16e-18 M=1
c2552 n95 n114 28.16e-18 M=1
c2553 n95 n108 56.24e-18 M=1
c2554 n95 n106 83.64e-18 M=1
c2555 n93 n202 88.64e-18 M=1
c2556 n93 n135 88.64e-18 M=1
c2557 n93 n125 88.64e-18 M=1
c2558 n88 n116 88.64e-18 M=1
c2559 n64 n215 55.84e-18 M=1
c2560 n61 n215 28.16e-18 M=1
c2561 n59 n201 28.16e-18 M=1
c2562 n59 n198 649.28e-18 M=1
c2563 n59 n190 55.84e-18 M=1
c2564 n59 n165 28.16e-18 M=1
c2565 n59 n159 28.16e-18 M=1
c2566 n59 n140 28.16e-18 M=1
c2567 n59 n133 28.16e-18 M=1
c2568 n59 n128 677.84e-18 M=1
c2569 n59 n116 725.44e-18 M=1
c2570 n59 n110 28.16e-18 M=1
c2571 n59 n104 28.16e-18 M=1
c2572 n59 n84 28.16e-18 M=1
c2573 n59 n78 28.16e-18 M=1
c2574 n57 n215 649.28e-18 M=1
c2575 n57 n202 88.64e-18 M=1
c2576 n57 n135 88.64e-18 M=1
c2577 n57 n125 88.64e-18 M=1
c2578 n57 n95 177.28e-18 M=1
c2579 n57 n93 88.64e-18 M=1
c2580 n57 n91 23.42e-18 M=1
c2581 n57 n72 191.7e-18 M=1
c2582 n53 n198 88.64e-18 M=1
c2583 n53 n168 88.64e-18 M=1
c2584 n53 n166 88.64e-18 M=1
c2585 n53 n150 28.16e-18 M=1
c2586 n53 n143 28.16e-18 M=1
c2587 n53 n136 56.64e-18 M=1
c2588 n53 n132 56.64e-18 M=1
c2589 n53 n128 233.92e-18 M=1
c2590 n53 n126 56.64e-18 M=1
c2591 n53 n119 56.64e-18 M=1
c2592 n53 n116 233.92e-18 M=1
c2593 n53 n112 28.16e-18 M=1
c2594 n53 n105 28.16e-18 M=1
c2595 n53 n88 88.64e-18 M=1
c2596 n53 n85 88.64e-18 M=1
c2597 n53 n59 408.32e-18 M=1
c2598 a9 n53 28.16e-18 M=1
c2599 a6 n202 28.16e-18 M=1
c2600 a5 n202 28.16e-18 M=1
c2601 a2 n358 28.16e-18 M=1
c2602 a1 n358 28.16e-18 M=1
c2603 b14 n209 28.16e-18 M=1
c2604 b13 n209 28.16e-18 M=1
c2605 b10 n53 28.16e-18 M=1
c2606 gnd n358 3.5306e-15 M=1
c2607 gnd n354 1.42658e-15 M=1
c2608 gnd n332 506.13e-18 M=1
c2609 gnd n330 466.48e-18 M=1
c2610 gnd n322 726.58e-18 M=1
c2611 gnd n291 4.19149e-15 M=1
c2612 gnd n284 2.54184e-15 M=1
c2613 gnd n281 2.54184e-15 M=1
c2614 gnd n272 4.19149e-15 M=1
c2615 gnd n251 726.58e-18 M=1
c2616 gnd n244 466.48e-18 M=1
c2617 gnd n241 506.13e-18 M=1
c2618 gnd n215 1.01008e-15 M=1
c2619 gnd n213 1.42658e-15 M=1
c2620 gnd n209 3.5306e-15 M=1
c2621 gnd n204 1.01008e-15 M=1
c2622 gnd n202 3.5306e-15 M=1
c2623 gnd n198 1.42658e-15 M=1
c2624 gnd n176 506.13e-18 M=1
c2625 gnd n174 466.48e-18 M=1
c2626 gnd n166 726.58e-18 M=1
c2627 gnd n135 4.19149e-15 M=1
c2628 gnd n128 2.54184e-15 M=1
c2629 gnd n125 2.54184e-15 M=1
c2630 gnd n116 4.19149e-15 M=1
c2631 gnd n95 726.58e-18 M=1
c2632 gnd n88 466.48e-18 M=1
c2633 gnd n85 506.13e-18 M=1
c2634 gnd n59 1.01008e-15 M=1
c2635 gnd n57 1.42658e-15 M=1
c2636 gnd n53 3.5306e-15 M=1
c2637 a14 n209 28.16e-18 M=1
c2638 a13 n209 28.16e-18 M=1
c2639 a10 n53 28.16e-18 M=1
c2640 cin n358 408.32e-18 M=1
c2641 cin n340 28.16e-18 M=1
c2642 cin n333 28.16e-18 M=1
c2643 cin n313 28.16e-18 M=1
c2644 cin n307 28.16e-18 M=1
c2645 cin n291 725.44e-18 M=1
c2646 cin n286 28.16e-18 M=1
c2647 cin n281 677.84e-18 M=1
c2648 cin n279 28.16e-18 M=1
c2649 cin n258 28.16e-18 M=1
c2650 cin n252 28.16e-18 M=1
c2651 cin n220 55.84e-18 M=1
c2652 cin n217 28.16e-18 M=1
c2653 cin n213 649.28e-18 M=1
c2654 cin s2 55.84e-18 M=1
c2655 cin s1 55.84e-18 M=1
c2656 cin s0 55.84e-18 M=1
c2657 cin gnd 1.01008e-15 M=1
c2658 s15 n204 55.84e-18 M=1
c2659 s14 n204 55.84e-18 M=1
c2660 s13 n204 55.84e-18 M=1
c2661 s12 n204 55.84e-18 M=1
c2662 s11 n59 55.84e-18 M=1
c2663 s10 n59 55.84e-18 M=1
c2664 b9 n53 28.16e-18 M=1
c2665 b6 n202 28.16e-18 M=1
c2666 b5 n202 28.16e-18 M=1
c2667 s9 n59 55.84e-18 M=1
c2668 s8 n59 55.84e-18 M=1
c2669 b2 n358 28.16e-18 M=1
c2670 s7 n215 55.84e-18 M=1
c2671 b1 n358 28.16e-18 M=1
c2672 s6 n215 55.84e-18 M=1
c2673 s5 n215 55.84e-18 M=1
c2674 s4 n215 55.84e-18 M=1
c2675 s3 cin 55.84e-18 M=1
c2676 s2 n401 42.88e-18 M=1
c2677 s2 n358 96.96e-18 M=1
c2678 s2 n298 105.825e-18 M=1
c2679 s2 n291 96.96e-18 M=1
c2680 s2 n285 42.88e-18 M=1
c2681 s2 n281 96.96e-18 M=1
c2682 s2 n279 42.88e-18 M=1
c2683 s2 n278 42.88e-18 M=1
c2684 s2 n270 106.455e-18 M=1
c2685 s2 n267 42.88e-18 M=1
c2686 s2 n251 96.96e-18 M=1
c2687 s1 n408 42.88e-18 M=1
c2688 s1 n407 42.88e-18 M=1
c2689 s1 n358 96.96e-18 M=1
c2690 s1 n317 42.88e-18 M=1
c2691 s1 n312 42.88e-18 M=1
c2692 s1 n311 42.88e-18 M=1
c2693 s1 n307 42.88e-18 M=1
c2694 s1 n305 42.88e-18 M=1
c2695 s1 n304 42.88e-18 M=1
c2696 s1 n298 84e-18 M=1
c2697 s1 n294 44.68e-18 M=1
c2698 s1 n291 205.32e-18 M=1
c2699 s0 n412 42.88e-18 M=1
c2700 s0 n358 96.96e-18 M=1
c2701 s0 n343 42.88e-18 M=1
c2702 s0 n337 160.765e-18 M=1
c2703 s0 n333 42.88e-18 M=1
c2704 s0 n330 96.96e-18 M=1
c2705 s0 n328 34.56e-18 M=1
c2706 s0 n325 55.9e-18 M=1
c2707 s0 n323 42.88e-18 M=1
c2708 a2 s2 79.84e-18 M=1
c2709 a1 s1 42.88e-18 M=1
c2710 gnd s2 353.32e-18 M=1
c2711 gnd s1 279.66e-18 M=1
c2712 gnd s0 411.04e-18 M=1
c2713 s15 n413 42.88e-18 M=1
c2714 s15 n354 96.96e-18 M=1
c2715 s15 n331 42.88e-18 M=1
c2716 s15 n327 87.68e-18 M=1
c2717 s15 n321 42.88e-18 M=1
c2718 s15 n318 42.88e-18 M=1
c2719 s15 n310 87.68e-18 M=1
c2720 s15 n284 96.96e-18 M=1
c2721 s15 n272 96.96e-18 M=1
c2722 s15 n209 96.96e-18 M=1
c2723 s15 gnd 434.3e-18 M=1
c2724 s14 n410 42.88e-18 M=1
c2725 s14 n322 96.96e-18 M=1
c2726 s14 n306 42.88e-18 M=1
c2727 s14 n303 106.455e-18 M=1
c2728 s14 n297 42.88e-18 M=1
c2729 s14 n296 42.88e-18 M=1
c2730 s14 n290 42.88e-18 M=1
c2731 s14 n284 96.96e-18 M=1
c2732 s14 n277 105.825e-18 M=1
c2733 s14 n272 96.96e-18 M=1
c2734 s14 n209 96.96e-18 M=1
c2735 s14 b14 42.88e-18 M=1
c2736 s14 gnd 353.32e-18 M=1
c2737 s14 a14 79.84e-18 M=1
c2738 s13 n403 42.88e-18 M=1
c2739 s13 n402 42.88e-18 M=1
c2740 s13 n277 84e-18 M=1
c2741 s13 n274 44.68e-18 M=1
c2742 s13 n272 205.32e-18 M=1
c2743 s13 n269 42.88e-18 M=1
c2744 s13 n268 42.88e-18 M=1
c2745 s13 n266 42.88e-18 M=1
c2746 s13 n263 42.88e-18 M=1
c2747 s13 n261 42.88e-18 M=1
c2748 s13 n256 42.88e-18 M=1
c2749 s13 n209 96.96e-18 M=1
c2750 s13 b13 127e-18 M=1
c2751 s13 gnd 279.66e-18 M=1
c2752 s13 a13 42.88e-18 M=1
c2753 s12 n398 42.88e-18 M=1
c2754 s12 n250 42.88e-18 M=1
c2755 s12 n246 34.56e-18 M=1
c2756 s12 n244 96.96e-18 M=1
c2757 s12 n243 55.9e-18 M=1
c2758 s12 n240 42.88e-18 M=1
c2759 s12 n236 160.765e-18 M=1
c2760 s12 n231 42.88e-18 M=1
c2761 s12 n209 96.96e-18 M=1
c2762 s12 gnd 408.58e-18 M=1
c2763 s11 n385 42.88e-18 M=1
c2764 s11 n198 96.96e-18 M=1
c2765 s11 n175 42.88e-18 M=1
c2766 s11 n171 87.68e-18 M=1
c2767 s11 n165 42.88e-18 M=1
c2768 s11 n162 42.88e-18 M=1
c2769 s11 n154 87.68e-18 M=1
c2770 s11 n128 96.96e-18 M=1
c2771 s11 n116 96.96e-18 M=1
c2772 s11 n53 96.96e-18 M=1
c2773 s11 gnd 434.3e-18 M=1
c2774 s10 n382 42.88e-18 M=1
c2775 s10 n166 96.96e-18 M=1
c2776 s10 n150 42.88e-18 M=1
c2777 s10 n147 106.455e-18 M=1
c2778 s10 n141 42.88e-18 M=1
c2779 s10 n140 42.88e-18 M=1
c2780 s10 n134 42.88e-18 M=1
c2781 s10 n128 96.96e-18 M=1
c2782 s10 n121 105.825e-18 M=1
c2783 s10 n116 96.96e-18 M=1
c2784 s10 n53 96.96e-18 M=1
c2785 s10 b10 42.88e-18 M=1
c2786 s10 gnd 353.32e-18 M=1
c2787 s10 a10 79.84e-18 M=1
c2788 s9 n375 42.88e-18 M=1
c2789 s9 n374 42.88e-18 M=1
c2790 s9 n121 84e-18 M=1
c2791 s9 n118 44.68e-18 M=1
c2792 s9 n116 205.32e-18 M=1
c2793 s9 n113 42.88e-18 M=1
c2794 s9 n112 42.88e-18 M=1
c2795 s9 n110 42.88e-18 M=1
c2796 s9 n107 42.88e-18 M=1
c2797 s9 n105 42.88e-18 M=1
c2798 s9 n100 42.88e-18 M=1
c2799 s9 n53 96.96e-18 M=1
c2800 s9 a9 42.88e-18 M=1
c2801 s9 gnd 279.66e-18 M=1
c2802 s9 b9 127e-18 M=1
c2803 s8 n370 42.88e-18 M=1
c2804 s8 n94 42.88e-18 M=1
c2805 s8 n90 34.56e-18 M=1
c2806 s8 n88 96.96e-18 M=1
c2807 s8 n87 55.9e-18 M=1
c2808 s8 n84 42.88e-18 M=1
c2809 s8 n80 160.765e-18 M=1
c2810 s8 n75 42.88e-18 M=1
c2811 s8 n53 96.96e-18 M=1
c2812 s8 gnd 408.58e-18 M=1
c2813 b2 s2 42.88e-18 M=1
c2814 s7 n369 42.88e-18 M=1
c2815 s7 n202 96.96e-18 M=1
c2816 s7 n135 96.96e-18 M=1
c2817 s7 n125 96.96e-18 M=1
c2818 s7 n108 87.68e-18 M=1
c2819 s7 n99 42.88e-18 M=1
c2820 s7 n96 42.88e-18 M=1
c2821 s7 n91 87.68e-18 M=1
c2822 s7 n86 42.88e-18 M=1
c2823 s7 n57 96.96e-18 M=1
c2824 s7 gnd 436.76e-18 M=1
c2825 b1 s1 127e-18 M=1
c2826 s6 n373 42.88e-18 M=1
c2827 s6 n202 96.96e-18 M=1
c2828 s6 n142 105.825e-18 M=1
c2829 s6 n135 96.96e-18 M=1
c2830 s6 n129 42.88e-18 M=1
c2831 s6 n125 96.96e-18 M=1
c2832 s6 n123 42.88e-18 M=1
c2833 s6 n122 42.88e-18 M=1
c2834 s6 n114 106.455e-18 M=1
c2835 s6 n111 42.88e-18 M=1
c2836 s6 n95 96.96e-18 M=1
c2837 s6 a6 79.84e-18 M=1
c2838 s6 gnd 355.78e-18 M=1
c2839 s6 b6 42.88e-18 M=1
c2840 s5 n380 42.88e-18 M=1
c2841 s5 n379 42.88e-18 M=1
c2842 s5 n202 96.96e-18 M=1
c2843 s5 n161 42.88e-18 M=1
c2844 s5 n156 42.88e-18 M=1
c2845 s5 n155 42.88e-18 M=1
c2846 s5 n151 42.88e-18 M=1
c2847 s5 n149 42.88e-18 M=1
c2848 s5 n148 42.88e-18 M=1
c2849 s5 n142 84e-18 M=1
c2850 s5 n138 44.68e-18 M=1
c2851 s5 n135 205.32e-18 M=1
c2852 s5 a5 42.88e-18 M=1
c2853 s5 gnd 282.12e-18 M=1
c2854 s5 b5 127e-18 M=1
c2855 vdd s2 356.91e-18 M=1
c2856 vdd s1 293.75e-18 M=1
c2857 vdd s0 386.935e-18 M=1
c2858 vdd s15 381.87e-18 M=1
c2859 vdd s14 356.91e-18 M=1
c2860 vdd s13 293.75e-18 M=1
c2861 vdd s12 386.935e-18 M=1
c2862 vdd s11 381.87e-18 M=1
c2863 vdd s10 356.91e-18 M=1
c2864 vdd s9 293.75e-18 M=1
c2865 vdd s8 386.935e-18 M=1
c2866 vdd s7 381.87e-18 M=1
c2867 vdd s6 356.91e-18 M=1
c2868 vdd s5 293.75e-18 M=1
c2869 s4 n384 42.88e-18 M=1
c2870 s4 n202 96.96e-18 M=1
c2871 s4 n187 42.88e-18 M=1
c2872 s4 n181 26.32e-18 M=1
c2873 s4 n177 42.88e-18 M=1
c2874 s4 n174 96.96e-18 M=1
c2875 s4 n172 34.56e-18 M=1
c2876 s4 n169 58.12e-18 M=1
c2877 s4 n167 42.88e-18 M=1
c2878 s4 gnd 498.86e-18 M=1
c2879 s4 vdd 442.685e-18 M=1
c2880 s3 n397 42.88e-18 M=1
c2881 s3 n358 96.96e-18 M=1
c2882 s3 n291 96.96e-18 M=1
c2883 s3 n281 96.96e-18 M=1
c2884 s3 n264 93.38e-18 M=1
c2885 s3 n255 42.88e-18 M=1
c2886 s3 n252 42.88e-18 M=1
c2887 s3 n247 93.38e-18 M=1
c2888 s3 n242 42.88e-18 M=1
c2889 s3 n213 96.96e-18 M=1
c2890 s3 gnd 446.28e-18 M=1
c2891 s3 vdd 393.86e-18 M=1
m2892 n54 n125 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2893 n55 n62 n53 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2894 n56 n57 n54 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2895 gnd n70 n55 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2896 n58 b8 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2897 n60 n68 n57 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2898 n53 a8 n58 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2899 gnd n73 n60 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2900 n63 a7 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2901 n57 b7 n63 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2902 n66 n74 n64 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2903 n67 n135 n65 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2904 gnd n76 n66 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2905 gnd n202 n67 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2906 n71 n215 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2907 n64 n61 n71 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2908 n72 n91 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2909 n76 n82 n72 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2910 n77 a8 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2911 n72 n99 n76 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2912 n79 b8 n77 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2913 n81 b7 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2914 n83 n96 s7 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2915 n86 a7 n81 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2916 gnd n102 n83 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2917 n89 n57 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2918 n90 n69 n87 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2919 n92 n59 s8 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2920 s7 n108 n89 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2921 n87 n80 n90 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2922 gnd n53 n92 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2923 gnd n75 n87 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2924 n97 n78 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2925 n98 a9 n94 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2926 s8 n84 n97 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2927 gnd b9 n98 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2928 n103 b6 n101 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2929 gnd a6 n103 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2930 n106 n122 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2931 n108 n114 n106 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2932 n106 n129 n108 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2933 n109 n123 s6 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2934 gnd n130 n109 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2935 n115 n125 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2936 n117 n90 s9 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2937 s6 n142 n115 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2938 n119 b9 n116 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2939 gnd n116 n117 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2940 n121 n100 n118 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2941 gnd a9 n119 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2942 n124 n104 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2943 n118 n113 n121 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2944 n126 n105 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2945 s9 n110 n124 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2946 n127 a6 n125 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2947 gnd n107 n118 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2948 n116 n112 n126 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2949 gnd b6 n127 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2950 n131 n111 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2951 n132 n143 n128 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2952 n125 n120 n131 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2953 gnd n150 n132 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2954 n136 b10 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2955 n137 n149 n135 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2956 n138 n155 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2957 n128 a10 n136 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2958 n139 n151 s5 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2959 gnd n156 n137 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2960 n142 n148 n138 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2961 gnd n157 n139 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2962 n144 a5 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2963 n138 n161 n142 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2964 n145 n135 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2965 n135 b5 n144 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2966 n146 n121 s10 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2967 s5 n172 n145 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2968 gnd n128 n146 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2969 n152 n133 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2970 s10 n140 n152 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2971 n154 n134 n153 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2972 n153 n147 n154 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2973 gnd n141 n153 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2974 n158 a10 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2975 n160 b10 n158 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2976 n163 b5 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2977 n164 n177 s4 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2978 n167 a5 n163 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2979 gnd n184 n164 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2980 n169 n187 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2981 n170 n202 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2982 n172 n181 n169 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2983 n173 n154 s11 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2984 s4 n215 n170 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2985 n169 n193 n172 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2986 gnd n198 n173 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2987 n178 n159 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2988 n180 a11 n175 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2989 s11 n165 n178 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2990 gnd b11 n180 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2991 n185 b4 n182 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2992 n186 n162 n183 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2993 gnd a4 n185 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2994 n183 n179 n186 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2995 gnd n171 n183 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m2996 n191 n201 n190 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2997 gnd n59 n191 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m2998 n195 n53 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m2999 n196 n186 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3000 n197 n116 n195 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3001 n190 n188 n196 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3002 n199 b11 n198 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3003 gnd a11 n199 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3004 n203 n189 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3005 n205 a4 n202 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3006 n198 n194 n203 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3007 gnd b4 n205 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3008 n207 n192 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3009 n208 n198 n206 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3010 n202 n200 n207 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3011 gnd n128 n208 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3012 n210 n281 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3013 n211 n218 n209 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3014 n212 n213 n210 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3015 gnd n226 n211 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3016 n214 b12 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3017 n216 n224 n213 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3018 n209 a12 n214 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3019 gnd n229 n216 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3020 n219 a3 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3021 n213 b3 n219 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3022 n222 n230 n220 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3023 n223 n291 n221 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3024 gnd n232 n222 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3025 gnd n358 n223 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3026 n227 cin gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3027 n220 n217 n227 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3028 n228 n247 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3029 n232 n238 n228 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3030 n233 a12 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3031 n228 n255 n232 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3032 n235 b12 n233 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3033 n237 b3 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3034 n239 n252 s3 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3035 n242 a3 n237 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3036 gnd n258 n239 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3037 n245 n213 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3038 n246 n225 n243 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3039 n248 n204 s12 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3040 s3 n264 n245 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3041 n243 n236 n246 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3042 gnd n209 n248 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3043 gnd n231 n243 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3044 n253 n234 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3045 n254 a13 n250 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3046 s12 n240 n253 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3047 gnd b13 n254 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3048 n259 b2 n257 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3049 gnd a2 n259 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3050 n262 n278 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3051 n264 n270 n262 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3052 n262 n285 n264 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3053 n265 n279 s2 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3054 gnd n286 n265 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3055 n271 n281 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3056 n273 n246 s13 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3057 s2 n298 n271 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3058 n275 b13 n272 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3059 gnd n272 n273 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3060 n277 n256 n274 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3061 gnd a13 n275 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3062 n280 n260 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3063 n274 n269 n277 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3064 n282 n261 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3065 s13 n266 n280 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3066 n283 a2 n281 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3067 gnd n263 n274 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3068 n272 n268 n282 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3069 gnd b2 n283 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3070 n287 n267 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3071 n288 n299 n284 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3072 n281 n276 n287 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3073 gnd n306 n288 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3074 n292 b14 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3075 n293 n305 n291 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3076 n294 n311 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3077 n284 a14 n292 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3078 n295 n307 s1 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3079 gnd n312 n293 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3080 n298 n304 n294 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3081 gnd n313 n295 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3082 n300 a1 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3083 n294 n317 n298 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3084 n301 n291 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3085 n291 b1 n300 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3086 n302 n277 s14 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3087 s1 n328 n301 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3088 gnd n284 n302 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3089 n308 n289 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3090 s14 n296 n308 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3091 n310 n290 n309 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3092 n309 n303 n310 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3093 gnd n297 n309 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3094 n314 a14 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3095 n316 b14 n314 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3096 n319 b1 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3097 n320 n333 s0 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3098 n323 a1 n319 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3099 gnd n340 n320 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3100 n325 n343 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3101 n326 n358 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3102 n328 n337 n325 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3103 n329 n310 s15 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3104 s0 cin n326 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3105 n325 n349 n328 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3106 gnd n354 n329 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3107 n334 n315 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3108 n336 a15 n331 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3109 s15 n321 n334 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3110 gnd b15 n336 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3111 n341 b0 n338 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3112 n342 n318 n339 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3113 gnd a0 n341 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3114 n339 n335 n342 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3115 gnd n327 n339 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3116 n347 n357 n346 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3117 gnd n204 n347 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3118 n351 n209 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3119 n352 n342 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3120 n353 n272 n351 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3121 n346 n344 n352 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3122 n355 b15 n354 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3123 gnd a15 n355 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3124 n359 n345 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3125 n360 a0 n358 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3126 n354 n350 n359 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3127 gnd b0 n360 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3128 n362 n348 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m3129 n363 n354 n361 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m3130 n358 n356 n362 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3131 gnd n284 n363 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m3132 gnd n64 n59 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3133 n61 n56 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=110e-15 AS=190e-15 PD=700e-9 PS=1.5e-6 M=1
m3134 gnd n65 n61 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=110e-15 PD=1.5e-6 PS=700e-9 M=1
m3135 gnd a8 n62 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3136 n69 n53 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3137 gnd b7 n68 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3138 gnd b8 n70 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3139 n75 n85 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3140 gnd a7 n73 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3141 gnd n61 n74 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3142 n78 n53 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3143 n80 n59 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3144 n84 n59 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3145 n85 n79 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3146 gnd n108 n82 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3147 gnd n94 n88 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3148 n93 n86 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3149 gnd n93 n91 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3150 gnd n101 n95 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3151 gnd n108 n96 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3152 gnd n57 n99 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3153 n100 n116 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3154 gnd n57 n102 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3155 n104 n116 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3156 n105 a9 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3157 n107 n88 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3158 n110 n90 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3159 n111 b6 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3160 n112 b9 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3161 n113 n90 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3162 gnd n142 n114 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3163 n120 a6 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3164 gnd n95 n122 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3165 gnd n142 n123 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3166 gnd n125 n129 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3167 gnd n125 n130 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3168 n133 n128 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3169 n134 n128 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3170 n140 n121 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3171 n141 n166 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3172 gnd a10 n143 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3173 n147 n121 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3174 gnd n172 n148 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3175 gnd b5 n149 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3176 gnd b10 n150 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3177 gnd n172 n151 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3178 gnd n174 n155 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3179 gnd a5 n156 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3180 gnd n135 n157 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3181 n159 n198 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3182 gnd n135 n161 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3183 n162 n198 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3184 n165 n154 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3185 n166 n160 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3186 n171 n168 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3187 gnd n175 n168 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3188 n174 n167 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3189 n179 n154 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3190 gnd n182 n176 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3191 gnd n215 n177 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3192 gnd n215 n181 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3193 gnd n202 n184 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3194 n188 n201 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3195 n189 a11 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3196 gnd n176 n187 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3197 n192 b4 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3198 n194 b11 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3199 gnd n202 n193 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3200 n200 a4 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3201 n201 n197 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=110e-15 AS=190e-15 PD=700e-9 PS=1.5e-6 M=1
m3202 gnd n206 n201 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=110e-15 PD=1.5e-6 PS=700e-9 M=1
m3203 n204 n190 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3204 gnd n220 n215 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3205 n217 n212 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=110e-15 AS=190e-15 PD=700e-9 PS=1.5e-6 M=1
m3206 gnd n221 n217 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=110e-15 PD=1.5e-6 PS=700e-9 M=1
m3207 gnd a12 n218 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3208 n225 n209 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3209 gnd b3 n224 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3210 gnd b12 n226 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3211 n231 n241 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3212 gnd a3 n229 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3213 gnd n217 n230 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3214 n234 n209 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3215 n236 n204 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3216 n240 n204 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3217 n241 n235 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3218 gnd n264 n238 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3219 gnd n250 n244 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3220 n249 n242 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3221 gnd n249 n247 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3222 gnd n257 n251 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3223 gnd n264 n252 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3224 gnd n213 n255 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3225 n256 n272 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3226 gnd n213 n258 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3227 n260 n272 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3228 n261 a13 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3229 n263 n244 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3230 n266 n246 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3231 n267 b2 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3232 n268 b13 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3233 n269 n246 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3234 gnd n298 n270 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3235 n276 a2 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3236 gnd n251 n278 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3237 gnd n298 n279 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3238 gnd n281 n285 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3239 gnd n281 n286 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3240 n289 n284 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3241 n290 n284 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3242 n296 n277 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3243 n297 n322 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3244 gnd a14 n299 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3245 n303 n277 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3246 gnd n328 n304 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3247 gnd b1 n305 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3248 gnd b14 n306 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3249 gnd n328 n307 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3250 gnd n330 n311 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3251 gnd a1 n312 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3252 gnd n291 n313 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3253 n315 n354 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3254 gnd n291 n317 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3255 n318 n354 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3256 n321 n310 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3257 n322 n316 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3258 n327 n324 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3259 gnd n331 n324 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3260 n330 n323 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3261 n335 n310 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3262 gnd n338 n332 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3263 gnd cin n333 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3264 gnd cin n337 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3265 gnd n358 n340 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3266 n344 n357 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3267 n345 a15 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3268 gnd n332 n343 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3269 n348 b0 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3270 n350 b15 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3271 gnd n358 n349 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3272 n356 a0 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3273 n357 n353 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=110e-15 AS=190e-15 PD=700e-9 PS=1.5e-6 M=1
m3274 gnd n361 n357 gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=110e-15 PD=1.5e-6 PS=700e-9 M=1
m3275 cout n346 gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m3276 vdd n62 n364 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3277 n364 n70 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3278 n53 b8 n364 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3279 vdd n68 n365 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3280 n364 a8 n53 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3281 n365 n73 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3282 n57 a7 n365 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3283 n365 b7 n57 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3284 vdd n74 n367 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3285 n367 n76 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3286 n64 n215 n367 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3287 n367 n61 n64 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3288 vdd n96 n369 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3289 n369 n102 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3290 s7 n57 n369 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3291 s8 n59 n370 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3292 n369 n108 s7 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3293 n370 n53 s8 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3294 vdd n78 n370 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3295 n370 n84 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3296 vdd n123 n373 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3297 n373 n130 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3298 s6 n125 n373 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3299 s9 n90 n374 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3300 n373 n142 s6 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3301 n116 b9 n375 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3302 n374 n116 s9 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3303 n375 a9 n116 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3304 vdd n104 n374 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3305 vdd n105 n375 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3306 n374 n110 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3307 n125 a6 n377 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3308 n375 n112 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3309 n377 b6 n125 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3310 vdd n111 n377 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3311 vdd n143 n378 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3312 n377 n120 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3313 n378 n150 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3314 n128 b10 n378 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3315 vdd n149 n379 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3316 n378 a10 n128 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3317 vdd n151 n380 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3318 n379 n156 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3319 n380 n157 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3320 n135 a5 n379 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3321 s5 n135 n380 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3322 n379 b5 n135 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3323 s10 n121 n382 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3324 n380 n172 s5 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3325 n382 n128 s10 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3326 vdd n133 n382 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3327 n382 n140 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3328 vdd n177 n384 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3329 n384 n184 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3330 s4 n202 n384 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3331 s11 n154 n385 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3332 n384 n215 s4 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3333 n385 n198 s11 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3334 vdd n159 n385 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3335 n385 n165 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3336 n190 n201 n388 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3337 n388 n59 n190 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3338 vdd n186 n388 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3339 n388 n188 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3340 n198 b11 n389 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3341 n389 a11 n198 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3342 vdd n189 n389 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3343 n202 a4 n391 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3344 n389 n194 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3345 n391 b4 n202 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3346 vdd n192 n391 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3347 n391 n200 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3348 vdd n218 n392 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3349 n392 n226 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3350 n209 b12 n392 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3351 vdd n224 n393 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3352 n392 a12 n209 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3353 n393 n229 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3354 n213 a3 n393 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3355 n393 b3 n213 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3356 vdd n230 n395 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3357 n395 n232 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3358 n220 cin n395 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3359 n395 n217 n220 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3360 vdd n252 n397 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3361 n397 n258 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3362 s3 n213 n397 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3363 s12 n204 n398 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3364 n397 n264 s3 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3365 n398 n209 s12 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3366 vdd n234 n398 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3367 n398 n240 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3368 vdd n279 n401 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3369 n401 n286 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3370 s2 n281 n401 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3371 s13 n246 n402 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3372 n401 n298 s2 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3373 n272 b13 n403 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3374 n402 n272 s13 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3375 n403 a13 n272 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3376 vdd n260 n402 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3377 vdd n261 n403 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3378 n402 n266 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3379 n281 a2 n405 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3380 n403 n268 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3381 n405 b2 n281 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3382 vdd n267 n405 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3383 vdd n299 n406 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3384 n405 n276 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3385 n406 n306 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3386 n284 b14 n406 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3387 vdd n305 n407 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3388 n406 a14 n284 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3389 vdd n307 n408 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3390 n407 n312 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3391 n408 n313 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3392 n291 a1 n407 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3393 s1 n291 n408 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3394 n407 b1 n291 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3395 s14 n277 n410 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3396 n408 n328 s1 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3397 n410 n284 s14 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3398 vdd n289 n410 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3399 n410 n296 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3400 vdd n333 n412 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3401 n412 n340 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3402 s0 n358 n412 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3403 s15 n310 n413 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3404 n412 cin s0 vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3405 n413 n354 s15 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3406 vdd n315 n413 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3407 n413 n321 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3408 n346 n357 n416 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3409 n416 n204 n346 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3410 vdd n342 n416 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3411 n416 n344 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3412 n354 b15 n417 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3413 n417 a15 n354 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3414 vdd n345 n417 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3415 n358 a0 n419 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m3416 n417 n350 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3417 n419 b0 n358 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3418 vdd n348 n419 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3419 n419 n356 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
m3420 vdd n64 n59 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3421 vdd a8 n62 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3422 n69 n53 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3423 vdd b7 n68 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3424 vdd b8 n70 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3425 n75 n85 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3426 vdd a7 n73 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3427 vdd n61 n74 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3428 n78 n53 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3429 n80 n59 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3430 n84 n59 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3431 n85 n79 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3432 vdd n108 n82 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3433 vdd n94 n88 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3434 n93 n86 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3435 vdd n93 n91 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3436 vdd n101 n95 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3437 vdd n108 n96 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3438 vdd n57 n99 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3439 n100 n116 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3440 vdd n57 n102 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3441 n104 n116 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3442 n105 a9 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3443 n107 n88 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3444 n110 n90 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3445 n111 b6 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3446 n112 b9 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3447 n113 n90 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3448 vdd n142 n114 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3449 n120 a6 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3450 vdd n95 n122 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3451 vdd n142 n123 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3452 vdd n125 n129 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3453 vdd n125 n130 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3454 n133 n128 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3455 n134 n128 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3456 n140 n121 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3457 n141 n166 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3458 vdd a10 n143 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3459 n147 n121 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3460 vdd n172 n148 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3461 vdd b5 n149 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3462 vdd b10 n150 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3463 vdd n172 n151 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3464 vdd n174 n155 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3465 vdd a5 n156 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3466 vdd n135 n157 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3467 n159 n198 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3468 vdd n135 n161 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3469 n162 n198 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3470 n165 n154 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3471 n166 n160 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3472 n171 n168 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3473 vdd n175 n168 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3474 n174 n167 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3475 n179 n154 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3476 vdd n182 n176 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3477 vdd n215 n177 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3478 vdd n215 n181 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3479 vdd n202 n184 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3480 n188 n201 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3481 n189 a11 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3482 vdd n176 n187 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3483 n192 b4 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3484 n194 b11 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3485 vdd n202 n193 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3486 n200 a4 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3487 n204 n190 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3488 vdd n220 n215 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3489 vdd a12 n218 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3490 n225 n209 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3491 vdd b3 n224 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3492 vdd b12 n226 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3493 n231 n241 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3494 vdd a3 n229 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3495 vdd n217 n230 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3496 n234 n209 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3497 n236 n204 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3498 n240 n204 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3499 n241 n235 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3500 vdd n264 n238 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3501 vdd n250 n244 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3502 n249 n242 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3503 vdd n249 n247 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3504 vdd n257 n251 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3505 vdd n264 n252 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3506 vdd n213 n255 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3507 n256 n272 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3508 vdd n213 n258 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3509 n260 n272 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3510 n261 a13 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3511 n263 n244 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3512 n266 n246 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3513 n267 b2 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3514 n268 b13 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3515 n269 n246 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3516 vdd n298 n270 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3517 n276 a2 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3518 vdd n251 n278 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3519 vdd n298 n279 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3520 vdd n281 n285 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3521 vdd n281 n286 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3522 n289 n284 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3523 n290 n284 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3524 n296 n277 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3525 n297 n322 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3526 vdd a14 n299 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3527 n303 n277 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3528 vdd n328 n304 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3529 vdd b1 n305 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3530 vdd b14 n306 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3531 vdd n328 n307 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3532 vdd n330 n311 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3533 vdd a1 n312 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3534 vdd n291 n313 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3535 n315 n354 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3536 vdd n291 n317 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3537 n318 n354 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3538 n321 n310 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3539 n322 n316 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3540 n327 n324 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3541 vdd n331 n324 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3542 n330 n323 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3543 n335 n310 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3544 vdd n338 n332 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3545 vdd cin n333 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3546 vdd cin n337 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3547 vdd n358 n340 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3548 n344 n357 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3549 n345 a15 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3550 vdd n332 n343 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3551 n348 b0 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3552 n350 b15 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3553 vdd n358 n349 vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3554 n356 a0 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3555 cout n346 vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m3556 n366 n56 vdd vdd tsmc20P L=200e-9 W=1.3e-6 AD=390e-15 AS=650e-15 PD=600e-9 PS=2.3e-6 M=1
m3557 n61 n65 n366 vdd tsmc20P L=200e-9 W=1.3e-6 AD=650e-15 AS=390e-15 PD=2.3e-6 PS=600e-9 M=1
m3558 n390 n197 n201 vdd tsmc20P L=200e-9 W=1.3e-6 AD=390e-15 AS=650e-15 PD=600e-9 PS=2.3e-6 M=1
m3559 vdd n206 n390 vdd tsmc20P L=200e-9 W=1.3e-6 AD=650e-15 AS=390e-15 PD=2.3e-6 PS=600e-9 M=1
m3560 n394 n212 vdd vdd tsmc20P L=200e-9 W=1.3e-6 AD=390e-15 AS=650e-15 PD=600e-9 PS=2.3e-6 M=1
m3561 n217 n221 n394 vdd tsmc20P L=200e-9 W=1.3e-6 AD=650e-15 AS=390e-15 PD=2.3e-6 PS=600e-9 M=1
m3562 n418 n353 n357 vdd tsmc20P L=200e-9 W=1.3e-6 AD=390e-15 AS=650e-15 PD=600e-9 PS=2.3e-6 M=1
m3563 vdd n361 n418 vdd tsmc20P L=200e-9 W=1.3e-6 AD=650e-15 AS=390e-15 PD=2.3e-6 PS=600e-9 M=1
m3564 vdd n91 n76 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3565 n368 n82 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3566 n76 n99 n368 vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3567 n371 n69 n90 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3568 vdd n80 n371 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3569 n90 n75 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3570 vdd n122 n108 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3571 n372 n114 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3572 n108 n129 n372 vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3573 n376 n100 n121 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3574 vdd n113 n376 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3575 n121 n107 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3576 vdd n155 n142 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3577 n381 n148 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3578 n142 n161 n381 vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3579 n383 n134 n154 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3580 vdd n147 n383 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3581 n154 n141 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3582 vdd n187 n172 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3583 n386 n181 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3584 n172 n193 n386 vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3585 n387 n162 n186 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3586 vdd n179 n387 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3587 n186 n171 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3588 vdd n247 n232 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3589 n396 n238 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3590 n232 n255 n396 vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3591 n399 n225 n246 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3592 vdd n236 n399 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3593 n246 n231 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3594 vdd n278 n264 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3595 n400 n270 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3596 n264 n285 n400 vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3597 n404 n256 n277 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3598 vdd n269 n404 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3599 n277 n263 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3600 vdd n311 n298 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3601 n409 n304 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3602 n298 n317 n409 vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3603 n411 n290 n310 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3604 vdd n303 n411 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3605 n310 n297 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3606 vdd n343 n328 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3607 n414 n337 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3608 n328 n349 n414 vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
m3609 n415 n318 n342 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m3610 vdd n335 n415 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m3611 n342 n327 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
.END
