** Generated for: hspiceD
** Generated on: Oct 17 23:26:19 2016
** Design library name: Assignment2
** Design cell name: q3_mux_sym_tb
** Design view name: schematic
.PARAM beta=1.764157


.TRAN 10e-9 3e-6 START=0.0

.OP

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20N.m"
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20P.m"

** Library name: Asst_6
** Cell name: q3_mux_schematic
** View name: schematic
.subckt q3_mux_schematic a b gnd f s vdd
mn2 f s_bar net24 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
mn0 f s net26 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
mn4 s_bar s gnd gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
mn3 net24 b gnd gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
mn1 net26 a gnd gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
mp3 net25 a vdd vdd tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
mp0 net23 b vdd vdd tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
mp2 f s_bar net25 vdd tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
mp1 f s net23 vdd tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
mp4 s_bar s vdd vdd tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
.ends q3_mux_schematic
** End of subcircuit definition.

** Library name: Assignment2
** Cell name: q3_mux_sym_tb
** View name: schematic
xi0 vdd b 0 net4 net1 vdd q3_mux_schematic
v1 vdd 0 DC=1.8
v0 net1 0 DC=0
c0 net4 0 5e-15 M=1
v2 b 0 PULSE 0 1.8 0 40e-9 40e-9 1e-6 2e-6
.END
