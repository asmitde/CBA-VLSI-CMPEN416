** Generated for: hspiceD
** Generated on: Nov 30 16:59:53 2016
** Design library name: Project_416
** Design cell name: full_adder
** Design view name: extracted


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20N.m"
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20P.m"

** Library name: Project_416
** Cell name: full_adder
** View name: extracted
m0 sum cin n17 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=400e-15 PD=600e-9 PS=1.8e-6 M=1
m1 n17 p sum vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m2 vdd n12 n17 vdd tsmc20P L=200e-9 W=800e-9 AD=240e-15 AS=240e-15 PD=600e-9 PS=600e-9 M=1
m3 n17 n13 vdd vdd tsmc20P L=200e-9 W=800e-9 AD=400e-15 AS=240e-15 PD=1.8e-6 PS=600e-9 M=1
c4 gnd n13 73.72e-18 M=1
c5 gnd n12 73.72e-18 M=1
c6 gnd n10 54.32e-18 M=1
c7 gnd n9 60.14e-18 M=1
c8 gnd n8 67.9e-18 M=1
c9 p gnd 124.16e-18 M=1
c10 g gnd 25.22e-18 M=1
c11 cin gnd 120.28e-18 M=1
c12 vdd n10 21.34e-18 M=1
c13 vdd p 62.08e-18 M=1
c14 vdd g 23.28e-18 M=1
c15 vdd cin 73.72e-18 M=1
c16 gnd n13 42.64e-18 M=1
c17 gnd n12 127e-18 M=1
c18 gnd n10 42.64e-18 M=1
c19 gnd n9 99.44e-18 M=1
c20 gnd n8 127.76e-18 M=1
c21 p gnd 225.68e-18 M=1
c22 g gnd 144.49e-18 M=1
c23 sum gnd 294.64e-18 M=1
c24 cin gnd 22.24e-18 M=1
c25 vdd n13 42.64e-18 M=1
c26 vdd n12 60.92e-18 M=1
c27 vdd n10 42.64e-18 M=1
c28 vdd n9 34.72e-18 M=1
c29 vdd n8 34.72e-18 M=1
c30 vdd gnd 528.83e-18 M=1
c31 vdd g 79.88e-18 M=1
c32 vdd sum 34.72e-18 M=1
c33 vdd cin 76.52e-18 M=1
c34 carry gnd 206.64e-18 M=1
c35 carry vdd 69.44e-18 M=1
c36 n13 n17 46.88e-18 M=1
c37 n12 n17 46.88e-18 M=1
c38 n12 n13 46.88e-18 M=1
c39 n10 n11 46.88e-18 M=1
c40 n9 n10 46.88e-18 M=1
c41 n8 n11 46.88e-18 M=1
c42 n8 n10 46.88e-18 M=1
c43 n8 n9 46.88e-18 M=1
c44 gnd n13 330.48e-18 M=1
c45 gnd n12 573.16e-18 M=1
c46 gnd n10 195e-18 M=1
c47 gnd n9 611.2e-18 M=1
c48 gnd n8 771.36e-18 M=1
c49 p n17 46.88e-18 M=1
c50 p n13 46.88e-18 M=1
c51 p n12 46.88e-18 M=1
c52 p gnd 3.66306e-15 M=1
c53 g n8 84.41e-18 M=1
c54 g gnd 502.1e-18 M=1
c55 g p 108.74e-18 M=1
c56 sum n17 85.36e-18 M=1
c57 sum n13 130.72e-18 M=1
c58 sum n12 130.72e-18 M=1
c59 sum gnd 2.3168e-15 M=1
c60 sum p 130.72e-18 M=1
c61 cin n17 46.88e-18 M=1
c62 cin n13 131.29e-18 M=1
c63 cin n12 131.29e-18 M=1
c64 cin n9 44.875e-18 M=1
c65 cin n8 44.875e-18 M=1
c66 cin gnd 2.65978e-15 M=1
c67 cin p 190.62e-18 M=1
c68 cin g 35e-18 M=1
c69 cin sum 46.88e-18 M=1
c70 vdd n17 85.36e-18 M=1
c71 vdd n13 59.44e-18 M=1
c72 vdd n12 35.88e-18 M=1
c73 vdd n10 199.32e-18 M=1
c74 vdd p 205.02e-18 M=1
c75 vdd g 261.33e-18 M=1
c76 vdd cin 1.34211e-15 M=1
c77 carry n11 85.36e-18 M=1
c78 carry n10 130.72e-18 M=1
c79 carry n9 130.72e-18 M=1
c80 carry n8 46.88e-18 M=1
c81 carry gnd 2.51635e-15 M=1
m82 carry n8 n11 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m83 n11 n10 carry gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m84 gnd n9 n11 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m85 n14 cin sum gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=300e-15 PD=600e-9 PS=1.6e-6 M=1
m86 gnd p n14 gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m87 n15 n12 gnd gnd tsmc20N L=200e-9 W=600e-9 AD=180e-15 AS=180e-15 PD=600e-9 PS=600e-9 M=1
m88 sum n13 n15 gnd tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=180e-15 PD=1.6e-6 PS=600e-9 M=1
m89 n8 p gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m90 n9 g gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m91 n10 cin gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m92 n12 p gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m93 n13 cin gnd gnd tsmc20N L=200e-9 W=300e-9 AD=190e-15 AS=190e-15 PD=1.5e-6 PS=1.5e-6 M=1
m94 n8 p vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m95 n9 g vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m96 n10 cin vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m97 n12 p vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m98 n13 cin vdd vdd tsmc20P L=200e-9 W=650e-9 AD=325e-15 AS=325e-15 PD=1.65e-6 PS=1.65e-6 M=1
m99 n16 n8 carry vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=375e-15 PD=600e-9 PS=1.75e-6 M=1
m100 vdd n10 n16 vdd tsmc20P L=200e-9 W=750e-9 AD=225e-15 AS=225e-15 PD=600e-9 PS=600e-9 M=1
m101 carry n9 vdd vdd tsmc20P L=200e-9 W=750e-9 AD=375e-15 AS=225e-15 PD=1.75e-6 PS=600e-9 M=1
.END
