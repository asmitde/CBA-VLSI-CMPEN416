** Generated for: hspiceD
** Generated on: Nov 23 20:50:49 2016
** Design library name: Project_416
** Design cell name: NAND2
** Design view name: schematic


.TRAN 10e-9 3e-6 START=0.0

.OP

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20N.m"
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20P.m"

** Library name: Project_416
** Cell name: NAND2
** View name: schematic
mn1 anandb a net14 gnd tsmc20N L=200e-9 W=600e-9 AD=150e-15 AS=150e-15 PD=1.6e-6 PS=1.6e-6 M=1
mn0 net14 b gnd gnd tsmc20N L=200e-9 W=600e-9 AD=150e-15 AS=150e-15 PD=1.6e-6 PS=1.6e-6 M=1
mp1 anandb b vdd vdd tsmc20P L=200e-9 W=950e-9 AD=475e-15 AS=475e-15 PD=2.9e-6 PS=2.9e-6 M=1
mp0 anandb a vdd vdd tsmc20P L=200e-9 W=950e-9 AD=475e-15 AS=475e-15 PD=2.9e-6 PS=2.9e-6 M=1
.END
