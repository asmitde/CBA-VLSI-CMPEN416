** Generated for: hspiceD
** Generated on: Sep 14 18:18:26 2016
** Design library name: Assignment2
** Design cell name: schema1
** Design view name: schematic
.GLOBAL vdd!


.PROBE DC
+    I1(m1)
.PROBE TRAN
+    I1(m1)
.DC v0 0.0 2.0 100e-3

.TRAN 200e-3 30.0 START=0.0

.OP

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20N.m"
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20P.m"

** Library name: Assignment2
** Cell name: schema1
** View name: schematic
m1 net6 net3 0 0 tsmc20N L=200e-9 W=300e-9 AD=150e-15 AS=150e-15 PD=1.6e-6 PS=1.6e-6 M=1
m0 net6 net3 net8 vdd! tsmc20P L=200e-9 W=300e-9 AD=150e-15 AS=150e-15 PD=1.6e-6 PS=1.6e-6 M=1
v0 net3 0 PULSE 0 1.8 0 1 1 3 6
v1 net8 0 DC=2
.END
