** Generated for: hspiceD
** Generated on: Nov 23 22:34:07 2016
** Design library name: Project_416
** Design cell name: NOR2_tb
** Design view name: schematic
.PARAM beta=3


.TRAN 10e-9 3e-6 START=0.0

.OP

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20N.m"
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20P.m"

** Library name: Project_416
** Cell name: NOR2
** View name: schematic
.subckt NOR2 a anorb b vdd gnd
m1 anorb b gnd gnd tsmc20N L=200e-9 W=300e-9 AD=150e-15 AS=150e-15 PD=1.6e-6 PS=1.6e-6 M=1
m0 anorb a gnd gnd tsmc20N L=200e-9 W=300e-9 AD=150e-15 AS=150e-15 PD=1.6e-6 PS=1.6e-6 M=1
mp1 net45 a vdd vdd tsmc20P L=200e-9 W=1.3e-6 AD=650e-15 AS=650e-15 PD=3.6e-6 PS=3.6e-6 M=1
mp0 anorb b net45 vdd tsmc20P L=200e-9 W=1.3e-6 AD=650e-15 AS=650e-15 PD=3.6e-6 PS=3.6e-6 M=1
.ends NOR2
** End of subcircuit definition.

** Library name: Project_416
** Cell name: NOR2_tb
** View name: schematic
xi0 net3 net5 net4 net2 0 NOR2
v1 net3 0 PULSE 1.8 0 0 40e-9 40e-9 1e-6 2e-6
v0 net4 0 PULSE 0 0 0 40e-9 40e-9 1e-6 2e-6
v2 net2 0 DC=1.8
c0 net5 0 5e-15 M=1
.END
