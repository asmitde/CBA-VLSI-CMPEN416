** Generated for: hspiceD
** Generated on: Oct 17 21:09:52 2016
** Design library name: Asst_5
** Design cell name: Asst5_Q2
** Design view name: schematic
.PARAM beta=3


.TRAN 10e-9 3e-6 START=0.0

.OP

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20N.m"
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20P.m"

** Library name: Asst_5
** Cell name: Asst5_Q2
** View name: schematic
mp4 s_bar s b b tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
mp3 net17 a b b tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
mp2 f s_bar net17 b tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
mp1 f s net15 b tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
mp0 net15 b b b tsmc20P L=200e-9 W='beta*600e-9' AD='((beta*600e-9)*2.5)*200e-9' AS='((beta*600e-9)*2.5)*200e-9' PD='(2*beta)*600e-9+1e-6' PS='(2*beta)*600e-9+1e-6' M=1
mn4 s_bar s 0 0 tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
mn3 net14 b 0 0 tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
mn2 f s_bar net14 0 tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
mn1 net16 a 0 0 tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
mn0 f s net16 0 tsmc20N L=200e-9 W=600e-9 AD=300e-15 AS=300e-15 PD=2.2e-6 PS=2.2e-6 M=1
v2 s 0 DC=1.8
vdd b 0 DC=1.8
c0 f 0 5e-15 M=1
v0 a 0 PULSE 1.8 0 0 40e-9 40e-9 1e-6 2e-6
.END
