** Generated for: hspiceD
** Generated on: Sep 14 22:55:08 2016
** Design library name: Assignment2
** Design cell name: Asst2_2
** Design view name: schematic
.PARAM vds=-1.8 vgs=0


.PROBE DC
+    I3(mp0)
.DC vds 0.0 -1.8 50e-3

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20N.m"
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20P.m"

** Library name: Assignment2
** Cell name: Asst2_2
** View name: schematic
mp0 0 net1 net2 0 tsmc20P L=200e-9 W=1e-6 AD=500e-15 AS=500e-15 PD=3e-6 PS=3e-6 M=1
v1 net1 0 DC=vgs
v0 net2 0 DC=vds
.END
