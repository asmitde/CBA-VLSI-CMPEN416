** Generated for: hspiceD
** Generated on: Sep 14 21:31:47 2016
** Design library name: Asst_2
** Design cell name: Asst_2_1
** Design view name: schematic
.PARAM vds=1.8 vgs=1.8


.PROBE DC
+    I1(mn0)
.DC vgs 0.0 1.8 50e-3

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20N.m"
.INCLUDE "/home/software/cadence-2009/local/ncsu-cdk-1.6.0.beta/models/hspice/public/tsmc20P.m"

** Library name: Asst_2
** Cell name: Asst_2_1
** View name: schematic
mn0 net02 net1 0 0 tsmc20N L=200e-9 W=1e-6 AD=500e-15 AS=500e-15 PD=3e-6 PS=3e-6 M=1
v1 net1 0 DC=vgs
v0 net02 0 DC=vds
.END
